-- Custom_qsys_vga_subsystem_char_buf_subsystem.vhd

-- Generated using ACDS version 18.1 646

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Custom_qsys_vga_subsystem_char_buf_subsystem is
	port (
		avalon_char_source_ready          : in  std_logic                     := '0';             --     avalon_char_source.ready
		avalon_char_source_startofpacket  : out std_logic;                                        --                       .startofpacket
		avalon_char_source_endofpacket    : out std_logic;                                        --                       .endofpacket
		avalon_char_source_valid          : out std_logic;                                        --                       .valid
		avalon_char_source_data           : out std_logic_vector(39 downto 0);                    --                       .data
		char_buf_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => '0'); -- char_buf_control_slave.address
		char_buf_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --                       .byteenable
		char_buf_control_slave_read       : in  std_logic                     := '0';             --                       .read
		char_buf_control_slave_write      : in  std_logic                     := '0';             --                       .write
		char_buf_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                       .writedata
		char_buf_control_slave_readdata   : out std_logic_vector(31 downto 0);                    --                       .readdata
		char_buf_slave_address            : in  std_logic_vector(10 downto 0) := (others => '0'); --         char_buf_slave.address
		char_buf_slave_clken              : in  std_logic                     := '0';             --                       .clken
		char_buf_slave_chipselect         : in  std_logic                     := '0';             --                       .chipselect
		char_buf_slave_write              : in  std_logic                     := '0';             --                       .write
		char_buf_slave_readdata           : out std_logic_vector(31 downto 0);                    --                       .readdata
		char_buf_slave_writedata          : in  std_logic_vector(31 downto 0) := (others => '0'); --                       .writedata
		char_buf_slave_byteenable         : in  std_logic_vector(3 downto 0)  := (others => '0'); --                       .byteenable
		sys_clk_clk                       : in  std_logic                     := '0';             --                sys_clk.clk
		sys_reset_reset_n                 : in  std_logic                     := '0'              --              sys_reset.reset_n
	);
end entity Custom_qsys_vga_subsystem_char_buf_subsystem;

architecture rtl of Custom_qsys_vga_subsystem_char_buf_subsystem is
	component Custom_qsys_vga_subsystem_char_buf_subsystem_onchip_memory2_0 is
		port (
			address     : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Custom_qsys_vga_subsystem_char_buf_subsystem_onchip_memory2_0;

	component Custom_qsys_vga_subsystem_char_buf_subsystem_video_ascii_to_image_0 is
		port (
			clk                     : in  std_logic                    := 'X';             -- clk
			reset                   : in  std_logic                    := 'X';             -- reset
			ascii_in_channel        : in  std_logic_vector(5 downto 0) := (others => 'X'); -- channel
			ascii_in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			ascii_in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			ascii_in_valid          : in  std_logic                    := 'X';             -- valid
			ascii_in_ready          : out std_logic;                                       -- ready
			ascii_in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			image_out_ready         : in  std_logic                    := 'X';             -- ready
			image_out_startofpacket : out std_logic;                                       -- startofpacket
			image_out_endofpacket   : out std_logic;                                       -- endofpacket
			image_out_valid         : out std_logic;                                       -- valid
			image_out_data          : out std_logic                                        -- data
		);
	end component Custom_qsys_vga_subsystem_char_buf_subsystem_video_ascii_to_image_0;

	component Custom_qsys_vga_subsystem_char_buf_subsystem_video_change_alpha_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(39 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(39 downto 0)                     -- data
		);
	end component Custom_qsys_vga_subsystem_char_buf_subsystem_video_change_alpha_0;

	component Custom_qsys_vga_subsystem_char_buf_subsystem_video_dma_controller_0 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(7 downto 0);                     -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component Custom_qsys_vga_subsystem_char_buf_subsystem_video_dma_controller_0;

	component Custom_qsys_vga_subsystem_char_buf_subsystem_video_rgb_resampler_0 is
		port (
			clk                      : in  std_logic                     := 'X'; -- clk
			reset                    : in  std_logic                     := 'X'; -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X'; -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X'; -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X'; -- valid
			stream_in_ready          : out std_logic;                            -- ready
			stream_in_data           : in  std_logic                     := 'X'; -- data
			slave_read               : in  std_logic                     := 'X'; -- read
			slave_readdata           : out std_logic_vector(31 downto 0);        -- readdata
			stream_out_ready         : in  std_logic                     := 'X'; -- ready
			stream_out_startofpacket : out std_logic;                            -- startofpacket
			stream_out_endofpacket   : out std_logic;                            -- endofpacket
			stream_out_valid         : out std_logic;                            -- valid
			stream_out_data          : out std_logic_vector(39 downto 0)         -- data
		);
	end component Custom_qsys_vga_subsystem_char_buf_subsystem_video_rgb_resampler_0;

	component Custom_qsys_vga_subsystem_char_buf_subsystem_video_scaler_0 is
		port (
			clk                      : in  std_logic                    := 'X';             -- clk
			reset                    : in  std_logic                    := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                    := 'X';             -- valid
			stream_in_ready          : out std_logic;                                       -- ready
			stream_in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                    := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                       -- startofpacket
			stream_out_endofpacket   : out std_logic;                                       -- endofpacket
			stream_out_valid         : out std_logic;                                       -- valid
			stream_out_data          : out std_logic_vector(7 downto 0);                    -- data
			stream_out_channel       : out std_logic_vector(5 downto 0)                     -- channel
		);
	end component Custom_qsys_vga_subsystem_char_buf_subsystem_video_scaler_0;

	component Custom_qsys_vga_subsystem_char_buf_subsystem_mm_interconnect_0 is
		port (
			sys_clk_clk_clk                                          : in  std_logic                     := 'X';             -- clk
			video_dma_controller_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			video_dma_controller_0_avalon_dma_master_address         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			video_dma_controller_0_avalon_dma_master_waitrequest     : out std_logic;                                        -- waitrequest
			video_dma_controller_0_avalon_dma_master_read            : in  std_logic                     := 'X';             -- read
			video_dma_controller_0_avalon_dma_master_readdata        : out std_logic_vector(7 downto 0);                     -- readdata
			video_dma_controller_0_avalon_dma_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			video_dma_controller_0_avalon_dma_master_lock            : in  std_logic                     := 'X';             -- lock
			onchip_memory2_0_s2_address                              : out std_logic_vector(10 downto 0);                    -- address
			onchip_memory2_0_s2_write                                : out std_logic;                                        -- write
			onchip_memory2_0_s2_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s2_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s2_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s2_chipselect                           : out std_logic;                                        -- chipselect
			onchip_memory2_0_s2_clken                                : out std_logic;                                        -- clken
			video_rgb_resampler_0_avalon_rgb_slave_read              : out std_logic;                                        -- read
			video_rgb_resampler_0_avalon_rgb_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Custom_qsys_vga_subsystem_char_buf_subsystem_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal video_ascii_to_image_0_avalon_image_source_valid                  : std_logic;                     -- video_ascii_to_image_0:image_out_valid -> video_rgb_resampler_0:stream_in_valid
	signal video_ascii_to_image_0_avalon_image_source_data                   : std_logic;                     -- video_ascii_to_image_0:image_out_data -> video_rgb_resampler_0:stream_in_data
	signal video_ascii_to_image_0_avalon_image_source_ready                  : std_logic;                     -- video_rgb_resampler_0:stream_in_ready -> video_ascii_to_image_0:image_out_ready
	signal video_ascii_to_image_0_avalon_image_source_startofpacket          : std_logic;                     -- video_ascii_to_image_0:image_out_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	signal video_ascii_to_image_0_avalon_image_source_endofpacket            : std_logic;                     -- video_ascii_to_image_0:image_out_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	signal video_dma_controller_0_avalon_pixel_source_valid                  : std_logic;                     -- video_dma_controller_0:stream_valid -> video_scaler_0:stream_in_valid
	signal video_dma_controller_0_avalon_pixel_source_data                   : std_logic_vector(7 downto 0);  -- video_dma_controller_0:stream_data -> video_scaler_0:stream_in_data
	signal video_dma_controller_0_avalon_pixel_source_ready                  : std_logic;                     -- video_scaler_0:stream_in_ready -> video_dma_controller_0:stream_ready
	signal video_dma_controller_0_avalon_pixel_source_startofpacket          : std_logic;                     -- video_dma_controller_0:stream_startofpacket -> video_scaler_0:stream_in_startofpacket
	signal video_dma_controller_0_avalon_pixel_source_endofpacket            : std_logic;                     -- video_dma_controller_0:stream_endofpacket -> video_scaler_0:stream_in_endofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_valid                     : std_logic;                     -- video_rgb_resampler_0:stream_out_valid -> video_change_alpha_0:stream_in_valid
	signal video_rgb_resampler_0_avalon_rgb_source_data                      : std_logic_vector(39 downto 0); -- video_rgb_resampler_0:stream_out_data -> video_change_alpha_0:stream_in_data
	signal video_rgb_resampler_0_avalon_rgb_source_ready                     : std_logic;                     -- video_change_alpha_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	signal video_rgb_resampler_0_avalon_rgb_source_startofpacket             : std_logic;                     -- video_rgb_resampler_0:stream_out_startofpacket -> video_change_alpha_0:stream_in_startofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_endofpacket               : std_logic;                     -- video_rgb_resampler_0:stream_out_endofpacket -> video_change_alpha_0:stream_in_endofpacket
	signal video_scaler_0_avalon_scaler_source_valid                         : std_logic;                     -- video_scaler_0:stream_out_valid -> video_ascii_to_image_0:ascii_in_valid
	signal video_scaler_0_avalon_scaler_source_data                          : std_logic_vector(7 downto 0);  -- video_scaler_0:stream_out_data -> video_ascii_to_image_0:ascii_in_data
	signal video_scaler_0_avalon_scaler_source_ready                         : std_logic;                     -- video_ascii_to_image_0:ascii_in_ready -> video_scaler_0:stream_out_ready
	signal video_scaler_0_avalon_scaler_source_channel                       : std_logic_vector(5 downto 0);  -- video_scaler_0:stream_out_channel -> video_ascii_to_image_0:ascii_in_channel
	signal video_scaler_0_avalon_scaler_source_startofpacket                 : std_logic;                     -- video_scaler_0:stream_out_startofpacket -> video_ascii_to_image_0:ascii_in_startofpacket
	signal video_scaler_0_avalon_scaler_source_endofpacket                   : std_logic;                     -- video_scaler_0:stream_out_endofpacket -> video_ascii_to_image_0:ascii_in_endofpacket
	signal video_dma_controller_0_avalon_dma_master_waitrequest              : std_logic;                     -- mm_interconnect_0:video_dma_controller_0_avalon_dma_master_waitrequest -> video_dma_controller_0:master_waitrequest
	signal video_dma_controller_0_avalon_dma_master_readdata                 : std_logic_vector(7 downto 0);  -- mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdata -> video_dma_controller_0:master_readdata
	signal video_dma_controller_0_avalon_dma_master_address                  : std_logic_vector(31 downto 0); -- video_dma_controller_0:master_address -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_address
	signal video_dma_controller_0_avalon_dma_master_read                     : std_logic;                     -- video_dma_controller_0:master_read -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_read
	signal video_dma_controller_0_avalon_dma_master_readdatavalid            : std_logic;                     -- mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdatavalid -> video_dma_controller_0:master_readdatavalid
	signal video_dma_controller_0_avalon_dma_master_lock                     : std_logic;                     -- video_dma_controller_0:master_arbiterlock -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_lock
	signal mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata : std_logic_vector(31 downto 0); -- video_rgb_resampler_0:slave_readdata -> mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_readdata
	signal mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read     : std_logic;                     -- mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_read -> video_rgb_resampler_0:slave_read
	signal mm_interconnect_0_onchip_memory2_0_s2_chipselect                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	signal mm_interconnect_0_onchip_memory2_0_s2_readdata                    : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	signal mm_interconnect_0_onchip_memory2_0_s2_address                     : std_logic_vector(10 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	signal mm_interconnect_0_onchip_memory2_0_s2_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	signal mm_interconnect_0_onchip_memory2_0_s2_write                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	signal mm_interconnect_0_onchip_memory2_0_s2_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	signal mm_interconnect_0_onchip_memory2_0_s2_clken                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:video_dma_controller_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset, video_ascii_to_image_0:reset, video_change_alpha_0:reset, video_dma_controller_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset]
	signal rst_controller_reset_out_reset_req                                : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal sys_reset_reset_n_ports_inv                                       : std_logic;                     -- sys_reset_reset_n:inv -> rst_controller:reset_in0

begin

	onchip_memory2_0 : component Custom_qsys_vga_subsystem_char_buf_subsystem_onchip_memory2_0
		port map (
			address     => char_buf_slave_address,                           --     s1.address
			clken       => char_buf_slave_clken,                             --       .clken
			chipselect  => char_buf_slave_chipselect,                        --       .chipselect
			write       => char_buf_slave_write,                             --       .write
			readdata    => char_buf_slave_readdata,                          --       .readdata
			writedata   => char_buf_slave_writedata,                         --       .writedata
			byteenable  => char_buf_slave_byteenable,                        --       .byteenable
			address2    => mm_interconnect_0_onchip_memory2_0_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_memory2_0_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_memory2_0_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_memory2_0_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_memory2_0_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_memory2_0_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_memory2_0_s2_byteenable, --       .byteenable
			clk         => sys_clk_clk,                                      --   clk1.clk
			reset       => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze      => '0'                                               -- (terminated)
		);

	video_ascii_to_image_0 : component Custom_qsys_vga_subsystem_char_buf_subsystem_video_ascii_to_image_0
		port map (
			clk                     => sys_clk_clk,                                              --                 clk.clk
			reset                   => rst_controller_reset_out_reset,                           --               reset.reset
			ascii_in_channel        => video_scaler_0_avalon_scaler_source_channel,              --   avalon_ascii_sink.channel
			ascii_in_startofpacket  => video_scaler_0_avalon_scaler_source_startofpacket,        --                    .startofpacket
			ascii_in_endofpacket    => video_scaler_0_avalon_scaler_source_endofpacket,          --                    .endofpacket
			ascii_in_valid          => video_scaler_0_avalon_scaler_source_valid,                --                    .valid
			ascii_in_ready          => video_scaler_0_avalon_scaler_source_ready,                --                    .ready
			ascii_in_data           => video_scaler_0_avalon_scaler_source_data,                 --                    .data
			image_out_ready         => video_ascii_to_image_0_avalon_image_source_ready,         -- avalon_image_source.ready
			image_out_startofpacket => video_ascii_to_image_0_avalon_image_source_startofpacket, --                    .startofpacket
			image_out_endofpacket   => video_ascii_to_image_0_avalon_image_source_endofpacket,   --                    .endofpacket
			image_out_valid         => video_ascii_to_image_0_avalon_image_source_valid,         --                    .valid
			image_out_data          => video_ascii_to_image_0_avalon_image_source_data           --                    .data
		);

	video_change_alpha_0 : component Custom_qsys_vga_subsystem_char_buf_subsystem_video_change_alpha_0
		port map (
			clk                      => sys_clk_clk,                                           --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                        --                     reset.reset
			stream_in_startofpacket  => video_rgb_resampler_0_avalon_rgb_source_startofpacket, --   avalon_apply_alpha_sink.startofpacket
			stream_in_endofpacket    => video_rgb_resampler_0_avalon_rgb_source_endofpacket,   --                          .endofpacket
			stream_in_valid          => video_rgb_resampler_0_avalon_rgb_source_valid,         --                          .valid
			stream_in_ready          => video_rgb_resampler_0_avalon_rgb_source_ready,         --                          .ready
			stream_in_data           => video_rgb_resampler_0_avalon_rgb_source_data,          --                          .data
			stream_out_ready         => avalon_char_source_ready,                              -- avalon_apply_alpha_source.ready
			stream_out_startofpacket => avalon_char_source_startofpacket,                      --                          .startofpacket
			stream_out_endofpacket   => avalon_char_source_endofpacket,                        --                          .endofpacket
			stream_out_valid         => avalon_char_source_valid,                              --                          .valid
			stream_out_data          => avalon_char_source_data                                --                          .data
		);

	video_dma_controller_0 : component Custom_qsys_vga_subsystem_char_buf_subsystem_video_dma_controller_0
		port map (
			clk                  => sys_clk_clk,                                              --                      clk.clk
			reset                => rst_controller_reset_out_reset,                           --                    reset.reset
			master_address       => video_dma_controller_0_avalon_dma_master_address,         --        avalon_dma_master.address
			master_waitrequest   => video_dma_controller_0_avalon_dma_master_waitrequest,     --                         .waitrequest
			master_arbiterlock   => video_dma_controller_0_avalon_dma_master_lock,            --                         .lock
			master_read          => video_dma_controller_0_avalon_dma_master_read,            --                         .read
			master_readdata      => video_dma_controller_0_avalon_dma_master_readdata,        --                         .readdata
			master_readdatavalid => video_dma_controller_0_avalon_dma_master_readdatavalid,   --                         .readdatavalid
			slave_address        => char_buf_control_slave_address,                           -- avalon_dma_control_slave.address
			slave_byteenable     => char_buf_control_slave_byteenable,                        --                         .byteenable
			slave_read           => char_buf_control_slave_read,                              --                         .read
			slave_write          => char_buf_control_slave_write,                             --                         .write
			slave_writedata      => char_buf_control_slave_writedata,                         --                         .writedata
			slave_readdata       => char_buf_control_slave_readdata,                          --                         .readdata
			stream_ready         => video_dma_controller_0_avalon_pixel_source_ready,         --      avalon_pixel_source.ready
			stream_data          => video_dma_controller_0_avalon_pixel_source_data,          --                         .data
			stream_startofpacket => video_dma_controller_0_avalon_pixel_source_startofpacket, --                         .startofpacket
			stream_endofpacket   => video_dma_controller_0_avalon_pixel_source_endofpacket,   --                         .endofpacket
			stream_valid         => video_dma_controller_0_avalon_pixel_source_valid          --                         .valid
		);

	video_rgb_resampler_0 : component Custom_qsys_vga_subsystem_char_buf_subsystem_video_rgb_resampler_0
		port map (
			clk                      => sys_clk_clk,                                                       --               clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --             reset.reset
			stream_in_startofpacket  => video_ascii_to_image_0_avalon_image_source_startofpacket,          --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => video_ascii_to_image_0_avalon_image_source_endofpacket,            --                  .endofpacket
			stream_in_valid          => video_ascii_to_image_0_avalon_image_source_valid,                  --                  .valid
			stream_in_ready          => video_ascii_to_image_0_avalon_image_source_ready,                  --                  .ready
			stream_in_data           => video_ascii_to_image_0_avalon_image_source_data,                   --                  .data
			slave_read               => mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read,     --  avalon_rgb_slave.read
			slave_readdata           => mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata, --                  .readdata
			stream_out_ready         => video_rgb_resampler_0_avalon_rgb_source_ready,                     -- avalon_rgb_source.ready
			stream_out_startofpacket => video_rgb_resampler_0_avalon_rgb_source_startofpacket,             --                  .startofpacket
			stream_out_endofpacket   => video_rgb_resampler_0_avalon_rgb_source_endofpacket,               --                  .endofpacket
			stream_out_valid         => video_rgb_resampler_0_avalon_rgb_source_valid,                     --                  .valid
			stream_out_data          => video_rgb_resampler_0_avalon_rgb_source_data                       --                  .data
		);

	video_scaler_0 : component Custom_qsys_vga_subsystem_char_buf_subsystem_video_scaler_0
		port map (
			clk                      => sys_clk_clk,                                              --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                           --                reset.reset
			stream_in_startofpacket  => video_dma_controller_0_avalon_pixel_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => video_dma_controller_0_avalon_pixel_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_dma_controller_0_avalon_pixel_source_valid,         --                     .valid
			stream_in_ready          => video_dma_controller_0_avalon_pixel_source_ready,         --                     .ready
			stream_in_data           => video_dma_controller_0_avalon_pixel_source_data,          --                     .data
			stream_out_ready         => video_scaler_0_avalon_scaler_source_ready,                -- avalon_scaler_source.ready
			stream_out_startofpacket => video_scaler_0_avalon_scaler_source_startofpacket,        --                     .startofpacket
			stream_out_endofpacket   => video_scaler_0_avalon_scaler_source_endofpacket,          --                     .endofpacket
			stream_out_valid         => video_scaler_0_avalon_scaler_source_valid,                --                     .valid
			stream_out_data          => video_scaler_0_avalon_scaler_source_data,                 --                     .data
			stream_out_channel       => video_scaler_0_avalon_scaler_source_channel               --                     .channel
		);

	mm_interconnect_0 : component Custom_qsys_vga_subsystem_char_buf_subsystem_mm_interconnect_0
		port map (
			sys_clk_clk_clk                                          => sys_clk_clk,                                                       --                                        sys_clk_clk.clk
			video_dma_controller_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                    -- video_dma_controller_0_reset_reset_bridge_in_reset.reset
			video_dma_controller_0_avalon_dma_master_address         => video_dma_controller_0_avalon_dma_master_address,                  --           video_dma_controller_0_avalon_dma_master.address
			video_dma_controller_0_avalon_dma_master_waitrequest     => video_dma_controller_0_avalon_dma_master_waitrequest,              --                                                   .waitrequest
			video_dma_controller_0_avalon_dma_master_read            => video_dma_controller_0_avalon_dma_master_read,                     --                                                   .read
			video_dma_controller_0_avalon_dma_master_readdata        => video_dma_controller_0_avalon_dma_master_readdata,                 --                                                   .readdata
			video_dma_controller_0_avalon_dma_master_readdatavalid   => video_dma_controller_0_avalon_dma_master_readdatavalid,            --                                                   .readdatavalid
			video_dma_controller_0_avalon_dma_master_lock            => video_dma_controller_0_avalon_dma_master_lock,                     --                                                   .lock
			onchip_memory2_0_s2_address                              => mm_interconnect_0_onchip_memory2_0_s2_address,                     --                                onchip_memory2_0_s2.address
			onchip_memory2_0_s2_write                                => mm_interconnect_0_onchip_memory2_0_s2_write,                       --                                                   .write
			onchip_memory2_0_s2_readdata                             => mm_interconnect_0_onchip_memory2_0_s2_readdata,                    --                                                   .readdata
			onchip_memory2_0_s2_writedata                            => mm_interconnect_0_onchip_memory2_0_s2_writedata,                   --                                                   .writedata
			onchip_memory2_0_s2_byteenable                           => mm_interconnect_0_onchip_memory2_0_s2_byteenable,                  --                                                   .byteenable
			onchip_memory2_0_s2_chipselect                           => mm_interconnect_0_onchip_memory2_0_s2_chipselect,                  --                                                   .chipselect
			onchip_memory2_0_s2_clken                                => mm_interconnect_0_onchip_memory2_0_s2_clken,                       --                                                   .clken
			video_rgb_resampler_0_avalon_rgb_slave_read              => mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read,     --             video_rgb_resampler_0_avalon_rgb_slave.read
			video_rgb_resampler_0_avalon_rgb_slave_readdata          => mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata  --                                                   .readdata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => sys_clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

end architecture rtl; -- of Custom_qsys_vga_subsystem_char_buf_subsystem
