library IEEE;
use IEEE.std_logic_1164.all;

entity HRV_buffer is
	port (clk, reset_n : in std_logic;
			HRV_in : in std_logic_vector(11 downto 0);
			HRV_out : out std_logic_vector(11 downto 0)
			);
end entity; 


architecture behavioural of HRV_buffer is
begin

	process (clk, reset_n)
		variable HRV_temp : std_logic_vector(11 downto 0);
	begin
	
		if reset_n = '0' then
			HRV_temp := (others => '0');
		
		elsif rising_edge(clk) then
		
			if HRV_in /= "000000000000" then
				HRV_temp := HRV_in;
			end if;
			
			HRV_out <= HRV_temp;
		end if;
	
	end process;

end architecture;