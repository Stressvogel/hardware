-- Custom_qsys.vhd

-- Generated using ACDS version 18.1 646

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Custom_qsys is
	port (
		hrv_hex0_readdata             : out   std_logic_vector(6 downto 0);                     --    hrv_hex0.readdata
		hrv_hex1_readdata             : out   std_logic_vector(6 downto 0);                     --    hrv_hex1.readdata
		hrv_hex2_readdata             : out   std_logic_vector(6 downto 0);                     --    hrv_hex2.readdata
		hrv_i2c_export                : inout std_logic_vector(1 downto 0)  := (others => '0'); --     hrv_i2c.export
		hrv_ledg_writeresponsevalid_n : out   std_logic;                                        --    hrv_ledg.writeresponsevalid_n
		hrv_ledr_readdata             : out   std_logic_vector(15 downto 0);                    --    hrv_ledr.readdata
		ps2_CLK                       : inout std_logic                     := '0';             --         ps2.CLK
		ps2_DAT                       : inout std_logic                     := '0';             --            .DAT
		pushbuttons_export            : in    std_logic_vector(3 downto 0)  := (others => '0'); -- pushbuttons.export
		ref_clk_clk                   : in    std_logic                     := '0';             --     ref_clk.clk
		ref_reset_reset               : in    std_logic                     := '0';             --   ref_reset.reset
		sdram_addr                    : out   std_logic_vector(12 downto 0);                    --       sdram.addr
		sdram_ba                      : out   std_logic_vector(1 downto 0);                     --            .ba
		sdram_cas_n                   : out   std_logic;                                        --            .cas_n
		sdram_cke                     : out   std_logic;                                        --            .cke
		sdram_cs_n                    : out   std_logic;                                        --            .cs_n
		sdram_dq                      : inout std_logic_vector(31 downto 0) := (others => '0'); --            .dq
		sdram_dqm                     : out   std_logic_vector(3 downto 0);                     --            .dqm
		sdram_ras_n                   : out   std_logic;                                        --            .ras_n
		sdram_we_n                    : out   std_logic;                                        --            .we_n
		sdram_clk_clk                 : out   std_logic;                                        --   sdram_clk.clk
		spi_MISO                      : in    std_logic                     := '0';             --         spi.MISO
		spi_MOSI                      : out   std_logic;                                        --            .MOSI
		spi_SCLK                      : out   std_logic;                                        --            .SCLK
		spi_SS_n                      : out   std_logic;                                        --            .SS_n
		spi_pio_export                : out   std_logic_vector(3 downto 0);                     --     spi_pio.export
		sram_DQ                       : inout std_logic_vector(15 downto 0) := (others => '0'); --        sram.DQ
		sram_ADDR                     : out   std_logic_vector(19 downto 0);                    --            .ADDR
		sram_LB_N                     : out   std_logic;                                        --            .LB_N
		sram_UB_N                     : out   std_logic;                                        --            .UB_N
		sram_CE_N                     : out   std_logic;                                        --            .CE_N
		sram_OE_N                     : out   std_logic;                                        --            .OE_N
		sram_WE_N                     : out   std_logic;                                        --            .WE_N
		vga_CLK                       : out   std_logic;                                        --         vga.CLK
		vga_HS                        : out   std_logic;                                        --            .HS
		vga_VS                        : out   std_logic;                                        --            .VS
		vga_BLANK                     : out   std_logic;                                        --            .BLANK
		vga_SYNC                      : out   std_logic;                                        --            .SYNC
		vga_R                         : out   std_logic_vector(7 downto 0);                     --            .R
		vga_G                         : out   std_logic_vector(7 downto 0);                     --            .G
		vga_B                         : out   std_logic_vector(7 downto 0)                      --            .B
	);
end entity Custom_qsys;

architecture rtl of Custom_qsys is
	component DE2_115 is
		port (
			csi_clock_clk              : in    std_logic                     := 'X';             -- clk
			csi_reset_reset            : in    std_logic                     := 'X';             -- reset
			avs_stress_level_address   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avs_stress_level_readdata  : out   std_logic_vector(15 downto 0);                    -- readdata
			avs_stress_level_write     : in    std_logic                     := 'X';             -- write
			avs_stress_level_writedata : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			I2C_GPIO                   : inout std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			HEX0_signal                : out   std_logic_vector(6 downto 0);                     -- readdata
			HEX1_signal                : out   std_logic_vector(6 downto 0);                     -- readdata
			HEX2_signal                : out   std_logic_vector(6 downto 0);                     -- readdata
			LEDG_signal                : out   std_logic;                                        -- writeresponsevalid_n
			LEDR_signal                : out   std_logic_vector(15 downto 0)                     -- readdata
		);
	end component DE2_115;

	component Custom_qsys_Interval_Timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Custom_qsys_Interval_Timer;

	component Custom_qsys_Interval_Timer_2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Custom_qsys_Interval_Timer_2;

	component Custom_qsys_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Custom_qsys_jtag_uart_0;

	component Custom_qsys_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(31 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Custom_qsys_nios2_gen2_0;

	component Custom_qsys_ps2_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic                     := 'X';             -- address
			chipselect  : in    std_logic                     := 'X';             -- chipselect
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			irq         : out   std_logic;                                        -- irq
			PS2_CLK     : inout std_logic                     := 'X';             -- export
			PS2_DAT     : inout std_logic                     := 'X'              -- export
		);
	end component Custom_qsys_ps2_0;

	component Custom_qsys_pushbuttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Custom_qsys_pushbuttons;

	component Custom_qsys_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component Custom_qsys_sdram_controller;

	component Custom_qsys_spi_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component Custom_qsys_spi_0;

	component Custom_qsys_spi_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component Custom_qsys_spi_pio;

	component Custom_qsys_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component Custom_qsys_sram_0;

	component Custom_qsys_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Custom_qsys_sys_sdram_pll_0;

	component Custom_qsys_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Custom_qsys_sysid_qsys_0;

	component Custom_qsys_vga_subsystem is
		port (
			bus_reset_reset_n                    : in  std_logic                     := 'X';             -- reset_n
			char_buffer_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			char_buffer_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			char_buffer_control_slave_read       : in  std_logic                     := 'X';             -- read
			char_buffer_control_slave_write      : in  std_logic                     := 'X';             -- write
			char_buffer_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			char_buffer_control_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			char_buffer_slave_address            : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			char_buffer_slave_clken              : in  std_logic                     := 'X';             -- clken
			char_buffer_slave_chipselect         : in  std_logic                     := 'X';             -- chipselect
			char_buffer_slave_write              : in  std_logic                     := 'X';             -- write
			char_buffer_slave_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			char_buffer_slave_writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			char_buffer_slave_byteenable         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			pixel_dma_control_slave_address      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pixel_dma_control_slave_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			pixel_dma_control_slave_read         : in  std_logic                     := 'X';             -- read
			pixel_dma_control_slave_write        : in  std_logic                     := 'X';             -- write
			pixel_dma_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pixel_dma_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			pixel_dma_master_address             : out std_logic_vector(31 downto 0);                    -- address
			pixel_dma_master_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			pixel_dma_master_lock                : out std_logic;                                        -- lock
			pixel_dma_master_read                : out std_logic;                                        -- read
			pixel_dma_master_readdata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			pixel_dma_master_readdatavalid       : in  std_logic                     := 'X';             -- readdatavalid
			rgb_slave_read                       : in  std_logic                     := 'X';             -- read
			rgb_slave_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			vga_CLK                              : out std_logic;                                        -- CLK
			vga_HS                               : out std_logic;                                        -- HS
			vga_VS                               : out std_logic;                                        -- VS
			vga_BLANK                            : out std_logic;                                        -- BLANK
			vga_SYNC                             : out std_logic;                                        -- SYNC
			vga_R                                : out std_logic_vector(7 downto 0);                     -- R
			vga_G                                : out std_logic_vector(7 downto 0);                     -- G
			vga_B                                : out std_logic_vector(7 downto 0);                     -- B
			vga_bus_clk_clk                      : in  std_logic                     := 'X';             -- clk
			vga_clk_clk                          : in  std_logic                     := 'X';             -- clk
			vga_reset_reset_n                    : in  std_logic                     := 'X'              -- reset_n
		);
	end component Custom_qsys_vga_subsystem;

	component Custom_qsys_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Custom_qsys_video_pll_0;

	component Custom_qsys_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk                         : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			ps2_0_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			vga_subsystem_bus_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                       : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                      : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address             : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest         : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			vga_subsystem_pixel_dma_master_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vga_subsystem_pixel_dma_master_waitrequest          : out std_logic;                                        -- waitrequest
			vga_subsystem_pixel_dma_master_read                 : in  std_logic                     := 'X';             -- read
			vga_subsystem_pixel_dma_master_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			vga_subsystem_pixel_dma_master_readdatavalid        : out std_logic;                                        -- readdatavalid
			vga_subsystem_pixel_dma_master_lock                 : in  std_logic                     := 'X';             -- lock
			Heartrate_Variability_stress_level_address          : out std_logic_vector(1 downto 0);                     -- address
			Heartrate_Variability_stress_level_write            : out std_logic;                                        -- write
			Heartrate_Variability_stress_level_readdata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Heartrate_Variability_stress_level_writedata        : out std_logic_vector(15 downto 0);                    -- writedata
			Interval_Timer_s1_address                           : out std_logic_vector(2 downto 0);                     -- address
			Interval_Timer_s1_write                             : out std_logic;                                        -- write
			Interval_Timer_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Interval_Timer_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			Interval_Timer_s1_chipselect                        : out std_logic;                                        -- chipselect
			Interval_Timer_2_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			Interval_Timer_2_s1_write                           : out std_logic;                                        -- write
			Interval_Timer_2_s1_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Interval_Timer_2_s1_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			Interval_Timer_2_s1_chipselect                      : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                 : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                  : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect            : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                  : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                   : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess            : out std_logic;                                        -- debugaccess
			ps2_0_avalon_ps2_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			ps2_0_avalon_ps2_slave_write                        : out std_logic;                                        -- write
			ps2_0_avalon_ps2_slave_read                         : out std_logic;                                        -- read
			ps2_0_avalon_ps2_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ps2_0_avalon_ps2_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			ps2_0_avalon_ps2_slave_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			ps2_0_avalon_ps2_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			ps2_0_avalon_ps2_slave_chipselect                   : out std_logic;                                        -- chipselect
			pushbuttons_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			pushbuttons_s1_write                                : out std_logic;                                        -- write
			pushbuttons_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pushbuttons_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			pushbuttons_s1_chipselect                           : out std_logic;                                        -- chipselect
			sdram_controller_s1_address                         : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                           : out std_logic;                                        -- write
			sdram_controller_s1_read                            : out std_logic;                                        -- read
			sdram_controller_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                   : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                      : out std_logic;                                        -- chipselect
			spi_0_spi_control_port_address                      : out std_logic_vector(2 downto 0);                     -- address
			spi_0_spi_control_port_write                        : out std_logic;                                        -- write
			spi_0_spi_control_port_read                         : out std_logic;                                        -- read
			spi_0_spi_control_port_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_0_spi_control_port_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			spi_0_spi_control_port_chipselect                   : out std_logic;                                        -- chipselect
			spi_pio_s1_address                                  : out std_logic_vector(2 downto 0);                     -- address
			spi_pio_s1_write                                    : out std_logic;                                        -- write
			spi_pio_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			spi_pio_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			spi_pio_s1_chipselect                               : out std_logic;                                        -- chipselect
			sram_0_avalon_sram_slave_address                    : out std_logic_vector(19 downto 0);                    -- address
			sram_0_avalon_sram_slave_write                      : out std_logic;                                        -- write
			sram_0_avalon_sram_slave_read                       : out std_logic;                                        -- read
			sram_0_avalon_sram_slave_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sram_0_avalon_sram_slave_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			sram_0_avalon_sram_slave_byteenable                 : out std_logic_vector(1 downto 0);                     -- byteenable
			sram_0_avalon_sram_slave_readdatavalid              : in  std_logic                     := 'X';             -- readdatavalid
			sysid_qsys_0_control_slave_address                  : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vga_subsystem_char_buffer_control_slave_address     : out std_logic_vector(1 downto 0);                     -- address
			vga_subsystem_char_buffer_control_slave_write       : out std_logic;                                        -- write
			vga_subsystem_char_buffer_control_slave_read        : out std_logic;                                        -- read
			vga_subsystem_char_buffer_control_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vga_subsystem_char_buffer_control_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			vga_subsystem_char_buffer_control_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			vga_subsystem_char_buffer_slave_address             : out std_logic_vector(10 downto 0);                    -- address
			vga_subsystem_char_buffer_slave_write               : out std_logic;                                        -- write
			vga_subsystem_char_buffer_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vga_subsystem_char_buffer_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			vga_subsystem_char_buffer_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			vga_subsystem_char_buffer_slave_chipselect          : out std_logic;                                        -- chipselect
			vga_subsystem_char_buffer_slave_clken               : out std_logic;                                        -- clken
			vga_subsystem_pixel_dma_control_slave_address       : out std_logic_vector(1 downto 0);                     -- address
			vga_subsystem_pixel_dma_control_slave_write         : out std_logic;                                        -- write
			vga_subsystem_pixel_dma_control_slave_read          : out std_logic;                                        -- read
			vga_subsystem_pixel_dma_control_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vga_subsystem_pixel_dma_control_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			vga_subsystem_pixel_dma_control_slave_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			vga_subsystem_rgb_slave_read                        : out std_logic;                                        -- read
			vga_subsystem_rgb_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Custom_qsys_mm_interconnect_0;

	component Custom_qsys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Custom_qsys_irq_mapper;

	component custom_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component custom_qsys_rst_controller;

	component custom_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component custom_qsys_rst_controller_001;

	signal sys_sdram_pll_0_sys_clk_clk                                          : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [Heartrate_Variability:csi_clock_clk, Interval_Timer:clk, Interval_Timer_2:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, nios2_gen2_0:clk, ps2_0:clk, pushbuttons:clk, rst_controller:clk, rst_controller_001:clk, sdram_controller:clk, spi_0:clk, spi_pio:clk, sram_0:clk, sysid_qsys_0:clock, vga_subsystem:vga_bus_clk_clk, video_pll_0:ref_clk_clk]
	signal video_pll_0_vga_clk_clk                                              : std_logic;                     -- video_pll_0:vga_clk_clk -> vga_subsystem:vga_clk_clk
	signal sys_sdram_pll_0_reset_source_reset                                   : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in0, sys_sdram_pll_0_reset_source_reset:in]
	signal video_pll_0_reset_source_reset                                       : std_logic;                     -- video_pll_0:reset_source_reset -> video_pll_0_reset_source_reset:in
	signal nios2_gen2_0_data_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                 : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                     : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                  : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                        : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                       : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                   : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                              : std_logic_vector(27 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                 : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal vga_subsystem_pixel_dma_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:vga_subsystem_pixel_dma_master_waitrequest -> vga_subsystem:pixel_dma_master_waitrequest
	signal vga_subsystem_pixel_dma_master_readdata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:vga_subsystem_pixel_dma_master_readdata -> vga_subsystem:pixel_dma_master_readdata
	signal vga_subsystem_pixel_dma_master_address                               : std_logic_vector(31 downto 0); -- vga_subsystem:pixel_dma_master_address -> mm_interconnect_0:vga_subsystem_pixel_dma_master_address
	signal vga_subsystem_pixel_dma_master_read                                  : std_logic;                     -- vga_subsystem:pixel_dma_master_read -> mm_interconnect_0:vga_subsystem_pixel_dma_master_read
	signal vga_subsystem_pixel_dma_master_readdatavalid                         : std_logic;                     -- mm_interconnect_0:vga_subsystem_pixel_dma_master_readdatavalid -> vga_subsystem:pixel_dma_master_readdatavalid
	signal vga_subsystem_pixel_dma_master_lock                                  : std_logic;                     -- vga_subsystem:pixel_dma_master_lock -> mm_interconnect_0:vga_subsystem_pixel_dma_master_lock
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata             : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest          : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                 : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_chipselect                  : std_logic;                     -- mm_interconnect_0:ps2_0_avalon_ps2_slave_chipselect -> ps2_0:chipselect
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_readdata                    : std_logic_vector(31 downto 0); -- ps2_0:readdata -> mm_interconnect_0:ps2_0_avalon_ps2_slave_readdata
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_waitrequest                 : std_logic;                     -- ps2_0:waitrequest -> mm_interconnect_0:ps2_0_avalon_ps2_slave_waitrequest
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_address                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ps2_0_avalon_ps2_slave_address -> ps2_0:address
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_read                        : std_logic;                     -- mm_interconnect_0:ps2_0_avalon_ps2_slave_read -> ps2_0:read
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ps2_0_avalon_ps2_slave_byteenable -> ps2_0:byteenable
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_write                       : std_logic;                     -- mm_interconnect_0:ps2_0_avalon_ps2_slave_write -> ps2_0:write
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:ps2_0_avalon_ps2_slave_writedata -> ps2_0:writedata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdata                  : std_logic_vector(15 downto 0); -- sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_address                   : std_logic_vector(19 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	signal mm_interconnect_0_sram_0_avalon_sram_slave_read                      : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	signal mm_interconnect_0_sram_0_avalon_sram_slave_byteenable                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid             : std_logic;                     -- sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	signal mm_interconnect_0_sram_0_avalon_sram_slave_write                     : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	signal mm_interconnect_0_sram_0_avalon_sram_slave_writedata                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	signal mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata   : std_logic_vector(31 downto 0); -- vga_subsystem:char_buffer_control_slave_readdata -> mm_interconnect_0:vga_subsystem_char_buffer_control_slave_readdata
	signal mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:vga_subsystem_char_buffer_control_slave_address -> vga_subsystem:char_buffer_control_slave_address
	signal mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read       : std_logic;                     -- mm_interconnect_0:vga_subsystem_char_buffer_control_slave_read -> vga_subsystem:char_buffer_control_slave_read
	signal mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:vga_subsystem_char_buffer_control_slave_byteenable -> vga_subsystem:char_buffer_control_slave_byteenable
	signal mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write      : std_logic;                     -- mm_interconnect_0:vga_subsystem_char_buffer_control_slave_write -> vga_subsystem:char_buffer_control_slave_write
	signal mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:vga_subsystem_char_buffer_control_slave_writedata -> vga_subsystem:char_buffer_control_slave_writedata
	signal mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect         : std_logic;                     -- mm_interconnect_0:vga_subsystem_char_buffer_slave_chipselect -> vga_subsystem:char_buffer_slave_chipselect
	signal mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata           : std_logic_vector(31 downto 0); -- vga_subsystem:char_buffer_slave_readdata -> mm_interconnect_0:vga_subsystem_char_buffer_slave_readdata
	signal mm_interconnect_0_vga_subsystem_char_buffer_slave_address            : std_logic_vector(10 downto 0); -- mm_interconnect_0:vga_subsystem_char_buffer_slave_address -> vga_subsystem:char_buffer_slave_address
	signal mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:vga_subsystem_char_buffer_slave_byteenable -> vga_subsystem:char_buffer_slave_byteenable
	signal mm_interconnect_0_vga_subsystem_char_buffer_slave_write              : std_logic;                     -- mm_interconnect_0:vga_subsystem_char_buffer_slave_write -> vga_subsystem:char_buffer_slave_write
	signal mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:vga_subsystem_char_buffer_slave_writedata -> vga_subsystem:char_buffer_slave_writedata
	signal mm_interconnect_0_vga_subsystem_char_buffer_slave_clken              : std_logic;                     -- mm_interconnect_0:vga_subsystem_char_buffer_slave_clken -> vga_subsystem:char_buffer_slave_clken
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata              : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest           : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess           : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                  : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata     : std_logic_vector(31 downto 0); -- vga_subsystem:pixel_dma_control_slave_readdata -> mm_interconnect_0:vga_subsystem_pixel_dma_control_slave_readdata
	signal mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:vga_subsystem_pixel_dma_control_slave_address -> vga_subsystem:pixel_dma_control_slave_address
	signal mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read         : std_logic;                     -- mm_interconnect_0:vga_subsystem_pixel_dma_control_slave_read -> vga_subsystem:pixel_dma_control_slave_read
	signal mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:vga_subsystem_pixel_dma_control_slave_byteenable -> vga_subsystem:pixel_dma_control_slave_byteenable
	signal mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write        : std_logic;                     -- mm_interconnect_0:vga_subsystem_pixel_dma_control_slave_write -> vga_subsystem:pixel_dma_control_slave_write
	signal mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:vga_subsystem_pixel_dma_control_slave_writedata -> vga_subsystem:pixel_dma_control_slave_writedata
	signal mm_interconnect_0_vga_subsystem_rgb_slave_readdata                   : std_logic_vector(31 downto 0); -- vga_subsystem:rgb_slave_readdata -> mm_interconnect_0:vga_subsystem_rgb_slave_readdata
	signal mm_interconnect_0_vga_subsystem_rgb_slave_read                       : std_logic;                     -- mm_interconnect_0:vga_subsystem_rgb_slave_read -> vga_subsystem:rgb_slave_read
	signal mm_interconnect_0_sdram_controller_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                       : std_logic_vector(31 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest                    : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                        : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                           : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid                  : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                          : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal mm_interconnect_0_spi_pio_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:spi_pio_s1_chipselect -> spi_pio:chipselect
	signal mm_interconnect_0_spi_pio_s1_readdata                                : std_logic_vector(31 downto 0); -- spi_pio:readdata -> mm_interconnect_0:spi_pio_s1_readdata
	signal mm_interconnect_0_spi_pio_s1_address                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_pio_s1_address -> spi_pio:address
	signal mm_interconnect_0_spi_pio_s1_write                                   : std_logic;                     -- mm_interconnect_0:spi_pio_s1_write -> mm_interconnect_0_spi_pio_s1_write:in
	signal mm_interconnect_0_spi_pio_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:spi_pio_s1_writedata -> spi_pio:writedata
	signal mm_interconnect_0_pushbuttons_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:pushbuttons_s1_chipselect -> pushbuttons:chipselect
	signal mm_interconnect_0_pushbuttons_s1_readdata                            : std_logic_vector(31 downto 0); -- pushbuttons:readdata -> mm_interconnect_0:pushbuttons_s1_readdata
	signal mm_interconnect_0_pushbuttons_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pushbuttons_s1_address -> pushbuttons:address
	signal mm_interconnect_0_pushbuttons_s1_write                               : std_logic;                     -- mm_interconnect_0:pushbuttons_s1_write -> mm_interconnect_0_pushbuttons_s1_write:in
	signal mm_interconnect_0_pushbuttons_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pushbuttons_s1_writedata -> pushbuttons:writedata
	signal mm_interconnect_0_interval_timer_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	signal mm_interconnect_0_interval_timer_s1_readdata                         : std_logic_vector(15 downto 0); -- Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	signal mm_interconnect_0_interval_timer_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	signal mm_interconnect_0_interval_timer_s1_write                            : std_logic;                     -- mm_interconnect_0:Interval_Timer_s1_write -> mm_interconnect_0_interval_timer_s1_write:in
	signal mm_interconnect_0_interval_timer_s1_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	signal mm_interconnect_0_interval_timer_2_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:Interval_Timer_2_s1_chipselect -> Interval_Timer_2:chipselect
	signal mm_interconnect_0_interval_timer_2_s1_readdata                       : std_logic_vector(15 downto 0); -- Interval_Timer_2:readdata -> mm_interconnect_0:Interval_Timer_2_s1_readdata
	signal mm_interconnect_0_interval_timer_2_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Interval_Timer_2_s1_address -> Interval_Timer_2:address
	signal mm_interconnect_0_interval_timer_2_s1_write                          : std_logic;                     -- mm_interconnect_0:Interval_Timer_2_s1_write -> mm_interconnect_0_interval_timer_2_s1_write:in
	signal mm_interconnect_0_interval_timer_2_s1_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:Interval_Timer_2_s1_writedata -> Interval_Timer_2:writedata
	signal mm_interconnect_0_spi_0_spi_control_port_chipselect                  : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	signal mm_interconnect_0_spi_0_spi_control_port_readdata                    : std_logic_vector(15 downto 0); -- spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	signal mm_interconnect_0_spi_0_spi_control_port_address                     : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	signal mm_interconnect_0_spi_0_spi_control_port_read                        : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_read -> mm_interconnect_0_spi_0_spi_control_port_read:in
	signal mm_interconnect_0_spi_0_spi_control_port_write                       : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_write -> mm_interconnect_0_spi_0_spi_control_port_write:in
	signal mm_interconnect_0_spi_0_spi_control_port_writedata                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	signal mm_interconnect_0_heartrate_variability_stress_level_readdata        : std_logic_vector(15 downto 0); -- Heartrate_Variability:avs_stress_level_readdata -> mm_interconnect_0:Heartrate_Variability_stress_level_readdata
	signal mm_interconnect_0_heartrate_variability_stress_level_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Heartrate_Variability_stress_level_address -> Heartrate_Variability:avs_stress_level_address
	signal mm_interconnect_0_heartrate_variability_stress_level_write           : std_logic;                     -- mm_interconnect_0:Heartrate_Variability_stress_level_write -> Heartrate_Variability:avs_stress_level_write
	signal mm_interconnect_0_heartrate_variability_stress_level_writedata       : std_logic_vector(15 downto 0); -- mm_interconnect_0:Heartrate_Variability_stress_level_writedata -> Heartrate_Variability:avs_stress_level_writedata
	signal irq_mapper_receiver0_irq                                             : std_logic;                     -- ps2_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                             : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                             : std_logic;                     -- spi_0:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                             : std_logic;                     -- pushbuttons:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                             : std_logic;                     -- Interval_Timer:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                             : std_logic;                     -- Interval_Timer_2:irq -> irq_mapper:receiver5_irq
	signal nios2_gen2_0_irq_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                       : std_logic;                     -- rst_controller:reset_out -> [Heartrate_Variability:csi_reset_reset, mm_interconnect_0:ps2_0_reset_reset_bridge_in_reset_reset, ps2_0:reset, rst_controller_reset_out_reset:in, sram_0:reset]
	signal nios2_gen2_0_debug_reset_request_reset                               : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in0
	signal rst_controller_001_reset_out_reset                                   : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:vga_subsystem_bus_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset, video_pll_0:ref_reset_reset]
	signal rst_controller_001_reset_out_reset_req                               : std_logic;                     -- rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal sys_sdram_pll_0_reset_source_reset_ports_inv                         : std_logic;                     -- sys_sdram_pll_0_reset_source_reset:inv -> vga_subsystem:bus_reset_reset_n
	signal video_pll_0_reset_source_reset_ports_inv                             : std_logic;                     -- video_pll_0_reset_source_reset:inv -> vga_subsystem:vga_reset_reset_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv                 : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv           : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal mm_interconnect_0_spi_pio_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_spi_pio_s1_write:inv -> spi_pio:write_n
	signal mm_interconnect_0_pushbuttons_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_pushbuttons_s1_write:inv -> pushbuttons:write_n
	signal mm_interconnect_0_interval_timer_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_interval_timer_s1_write:inv -> Interval_Timer:write_n
	signal mm_interconnect_0_interval_timer_2_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_interval_timer_2_s1_write:inv -> Interval_Timer_2:write_n
	signal mm_interconnect_0_spi_0_spi_control_port_read_ports_inv              : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_read:inv -> spi_0:read_n
	signal mm_interconnect_0_spi_0_spi_control_port_write_ports_inv             : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_write:inv -> spi_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                             : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Interval_Timer:reset_n, pushbuttons:reset_n, sdram_controller:reset_n, spi_0:reset_n, spi_pio:reset_n, sysid_qsys_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                         : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [Interval_Timer_2:reset_n, jtag_uart_0:rst_n, nios2_gen2_0:reset_n]

begin

	heartrate_variability : component DE2_115
		port map (
			csi_clock_clk              => sys_sdram_pll_0_sys_clk_clk,                                    --        clock.clk
			csi_reset_reset            => rst_controller_reset_out_reset,                                 --  reset_reset.reset
			avs_stress_level_address   => mm_interconnect_0_heartrate_variability_stress_level_address,   -- stress_level.address
			avs_stress_level_readdata  => mm_interconnect_0_heartrate_variability_stress_level_readdata,  --             .readdata
			avs_stress_level_write     => mm_interconnect_0_heartrate_variability_stress_level_write,     --             .write
			avs_stress_level_writedata => mm_interconnect_0_heartrate_variability_stress_level_writedata, --             .writedata
			I2C_GPIO                   => hrv_i2c_export,                                                 --          I2C.export
			HEX0_signal                => hrv_hex0_readdata,                                              --         HEX0.readdata
			HEX1_signal                => hrv_hex1_readdata,                                              --         HEX1.readdata
			HEX2_signal                => hrv_hex2_readdata,                                              --         HEX2.readdata
			LEDG_signal                => hrv_ledg_writeresponsevalid_n,                                  --         LEDG.writeresponsevalid_n
			LEDR_signal                => hrv_ledr_readdata                                               --         LEDR.readdata
		);

	interval_timer : component Custom_qsys_Interval_Timer
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                         --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_0_interval_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_interval_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_interval_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_interval_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_interval_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                             --   irq.irq
		);

	interval_timer_2 : component Custom_qsys_Interval_Timer_2
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                           --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,          -- reset.reset_n
			address    => mm_interconnect_0_interval_timer_2_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_interval_timer_2_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_interval_timer_2_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_interval_timer_2_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_interval_timer_2_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                               --   irq.irq
		);

	jtag_uart_0 : component Custom_qsys_jtag_uart_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                     --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component Custom_qsys_nios2_gen2_0
		port map (
			clk                                 => sys_sdram_pll_0_sys_clk_clk,                                --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	ps2_0 : component Custom_qsys_ps2_0
		port map (
			clk         => sys_sdram_pll_0_sys_clk_clk,                          --                clk.clk
			reset       => rst_controller_reset_out_reset,                       --              reset.reset
			address     => mm_interconnect_0_ps2_0_avalon_ps2_slave_address(0),  --   avalon_ps2_slave.address
			chipselect  => mm_interconnect_0_ps2_0_avalon_ps2_slave_chipselect,  --                   .chipselect
			byteenable  => mm_interconnect_0_ps2_0_avalon_ps2_slave_byteenable,  --                   .byteenable
			read        => mm_interconnect_0_ps2_0_avalon_ps2_slave_read,        --                   .read
			write       => mm_interconnect_0_ps2_0_avalon_ps2_slave_write,       --                   .write
			writedata   => mm_interconnect_0_ps2_0_avalon_ps2_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_ps2_0_avalon_ps2_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_ps2_0_avalon_ps2_slave_waitrequest, --                   .waitrequest
			irq         => irq_mapper_receiver0_irq,                             --          interrupt.irq
			PS2_CLK     => ps2_CLK,                                              -- external_interface.export
			PS2_DAT     => ps2_DAT                                               --                   .export
		);

	pushbuttons : component Custom_qsys_pushbuttons
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_pushbuttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pushbuttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pushbuttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pushbuttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pushbuttons_s1_readdata,        --                    .readdata
			in_port    => pushbuttons_export,                               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                          --                 irq.irq
		);

	sdram_controller : component Custom_qsys_sdram_controller
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                                 --  wire.export
			zs_ba          => sdram_ba,                                                   --      .export
			zs_cas_n       => sdram_cas_n,                                                --      .export
			zs_cke         => sdram_cke,                                                  --      .export
			zs_cs_n        => sdram_cs_n,                                                 --      .export
			zs_dq          => sdram_dq,                                                   --      .export
			zs_dqm         => sdram_dqm,                                                  --      .export
			zs_ras_n       => sdram_ras_n,                                                --      .export
			zs_we_n        => sdram_we_n                                                  --      .export
		);

	spi_0 : component Custom_qsys_spi_0
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,                              --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                 --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_0_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_0_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_0_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_0_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_0_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_0_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver2_irq,                                 --              irq.irq
			MISO          => spi_MISO,                                                 --         external.export
			MOSI          => spi_MOSI,                                                 --                 .export
			SCLK          => spi_SCLK,                                                 --                 .export
			SS_n          => spi_SS_n                                                  --                 .export
		);

	spi_pio : component Custom_qsys_spi_pio
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_spi_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_spi_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_spi_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_spi_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_spi_pio_s1_readdata,        --                    .readdata
			out_port   => spi_pio_export                                -- external_connection.export
		);

	sram_0 : component Custom_qsys_sram_0
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,                              --                clk.clk
			reset         => rst_controller_reset_out_reset,                           --              reset.reset
			SRAM_DQ       => sram_DQ,                                                  -- external_interface.export
			SRAM_ADDR     => sram_ADDR,                                                --                   .export
			SRAM_LB_N     => sram_LB_N,                                                --                   .export
			SRAM_UB_N     => sram_UB_N,                                                --                   .export
			SRAM_CE_N     => sram_CE_N,                                                --                   .export
			SRAM_OE_N     => sram_OE_N,                                                --                   .export
			SRAM_WE_N     => sram_WE_N,                                                --                   .export
			address       => mm_interconnect_0_sram_0_avalon_sram_slave_address,       --  avalon_sram_slave.address
			byteenable    => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,    --                   .byteenable
			read          => mm_interconnect_0_sram_0_avalon_sram_slave_read,          --                   .read
			write         => mm_interconnect_0_sram_0_avalon_sram_slave_write,         --                   .write
			writedata     => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,     --                   .writedata
			readdata      => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,      --                   .readdata
			readdatavalid => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid  --                   .readdatavalid
		);

	sys_sdram_pll_0 : component Custom_qsys_sys_sdram_pll_0
		port map (
			ref_clk_clk        => ref_clk_clk,                        --      ref_clk.clk
			ref_reset_reset    => ref_reset_reset,                    --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	sysid_qsys_0 : component Custom_qsys_sysid_qsys_0
		port map (
			clock    => sys_sdram_pll_0_sys_clk_clk,                             --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	vga_subsystem : component Custom_qsys_vga_subsystem
		port map (
			bus_reset_reset_n                    => sys_sdram_pll_0_reset_source_reset_ports_inv,                         --                 bus_reset.reset_n
			char_buffer_control_slave_address    => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address,    -- char_buffer_control_slave.address
			char_buffer_control_slave_byteenable => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable, --                          .byteenable
			char_buffer_control_slave_read       => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read,       --                          .read
			char_buffer_control_slave_write      => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write,      --                          .write
			char_buffer_control_slave_writedata  => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata,  --                          .writedata
			char_buffer_control_slave_readdata   => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata,   --                          .readdata
			char_buffer_slave_address            => mm_interconnect_0_vga_subsystem_char_buffer_slave_address,            --         char_buffer_slave.address
			char_buffer_slave_clken              => mm_interconnect_0_vga_subsystem_char_buffer_slave_clken,              --                          .clken
			char_buffer_slave_chipselect         => mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect,         --                          .chipselect
			char_buffer_slave_write              => mm_interconnect_0_vga_subsystem_char_buffer_slave_write,              --                          .write
			char_buffer_slave_readdata           => mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata,           --                          .readdata
			char_buffer_slave_writedata          => mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata,          --                          .writedata
			char_buffer_slave_byteenable         => mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable,         --                          .byteenable
			pixel_dma_control_slave_address      => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address,      --   pixel_dma_control_slave.address
			pixel_dma_control_slave_byteenable   => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable,   --                          .byteenable
			pixel_dma_control_slave_read         => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read,         --                          .read
			pixel_dma_control_slave_write        => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write,        --                          .write
			pixel_dma_control_slave_writedata    => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata,    --                          .writedata
			pixel_dma_control_slave_readdata     => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata,     --                          .readdata
			pixel_dma_master_address             => vga_subsystem_pixel_dma_master_address,                               --          pixel_dma_master.address
			pixel_dma_master_waitrequest         => vga_subsystem_pixel_dma_master_waitrequest,                           --                          .waitrequest
			pixel_dma_master_lock                => vga_subsystem_pixel_dma_master_lock,                                  --                          .lock
			pixel_dma_master_read                => vga_subsystem_pixel_dma_master_read,                                  --                          .read
			pixel_dma_master_readdata            => vga_subsystem_pixel_dma_master_readdata,                              --                          .readdata
			pixel_dma_master_readdatavalid       => vga_subsystem_pixel_dma_master_readdatavalid,                         --                          .readdatavalid
			rgb_slave_read                       => mm_interconnect_0_vga_subsystem_rgb_slave_read,                       --                 rgb_slave.read
			rgb_slave_readdata                   => mm_interconnect_0_vga_subsystem_rgb_slave_readdata,                   --                          .readdata
			vga_CLK                              => vga_CLK,                                                              --                       vga.CLK
			vga_HS                               => vga_HS,                                                               --                          .HS
			vga_VS                               => vga_VS,                                                               --                          .VS
			vga_BLANK                            => vga_BLANK,                                                            --                          .BLANK
			vga_SYNC                             => vga_SYNC,                                                             --                          .SYNC
			vga_R                                => vga_R,                                                                --                          .R
			vga_G                                => vga_G,                                                                --                          .G
			vga_B                                => vga_B,                                                                --                          .B
			vga_bus_clk_clk                      => sys_sdram_pll_0_sys_clk_clk,                                          --               vga_bus_clk.clk
			vga_clk_clk                          => video_pll_0_vga_clk_clk,                                              --                   vga_clk.clk
			vga_reset_reset_n                    => video_pll_0_reset_source_reset_ports_inv                              --                 vga_reset.reset_n
		);

	video_pll_0 : component Custom_qsys_video_pll_0
		port map (
			ref_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => rst_controller_001_reset_out_reset, --    ref_reset.reset
			vga_clk_clk        => video_pll_0_vga_clk_clk,            --      vga_clk.clk
			reset_source_reset => video_pll_0_reset_source_reset      -- reset_source.reset
		);

	mm_interconnect_0 : component Custom_qsys_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk                         => sys_sdram_pll_0_sys_clk_clk,                                          --                       sys_sdram_pll_0_sys_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset      => rst_controller_001_reset_out_reset,                                   --      nios2_gen2_0_reset_reset_bridge_in_reset.reset
			ps2_0_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                                       --             ps2_0_reset_reset_bridge_in_reset.reset
			vga_subsystem_bus_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                   -- vga_subsystem_bus_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                    => nios2_gen2_0_data_master_address,                                     --                      nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                => nios2_gen2_0_data_master_waitrequest,                                 --                                              .waitrequest
			nios2_gen2_0_data_master_byteenable                 => nios2_gen2_0_data_master_byteenable,                                  --                                              .byteenable
			nios2_gen2_0_data_master_read                       => nios2_gen2_0_data_master_read,                                        --                                              .read
			nios2_gen2_0_data_master_readdata                   => nios2_gen2_0_data_master_readdata,                                    --                                              .readdata
			nios2_gen2_0_data_master_write                      => nios2_gen2_0_data_master_write,                                       --                                              .write
			nios2_gen2_0_data_master_writedata                  => nios2_gen2_0_data_master_writedata,                                   --                                              .writedata
			nios2_gen2_0_data_master_debugaccess                => nios2_gen2_0_data_master_debugaccess,                                 --                                              .debugaccess
			nios2_gen2_0_instruction_master_address             => nios2_gen2_0_instruction_master_address,                              --               nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest         => nios2_gen2_0_instruction_master_waitrequest,                          --                                              .waitrequest
			nios2_gen2_0_instruction_master_read                => nios2_gen2_0_instruction_master_read,                                 --                                              .read
			nios2_gen2_0_instruction_master_readdata            => nios2_gen2_0_instruction_master_readdata,                             --                                              .readdata
			vga_subsystem_pixel_dma_master_address              => vga_subsystem_pixel_dma_master_address,                               --                vga_subsystem_pixel_dma_master.address
			vga_subsystem_pixel_dma_master_waitrequest          => vga_subsystem_pixel_dma_master_waitrequest,                           --                                              .waitrequest
			vga_subsystem_pixel_dma_master_read                 => vga_subsystem_pixel_dma_master_read,                                  --                                              .read
			vga_subsystem_pixel_dma_master_readdata             => vga_subsystem_pixel_dma_master_readdata,                              --                                              .readdata
			vga_subsystem_pixel_dma_master_readdatavalid        => vga_subsystem_pixel_dma_master_readdatavalid,                         --                                              .readdatavalid
			vga_subsystem_pixel_dma_master_lock                 => vga_subsystem_pixel_dma_master_lock,                                  --                                              .lock
			Heartrate_Variability_stress_level_address          => mm_interconnect_0_heartrate_variability_stress_level_address,         --            Heartrate_Variability_stress_level.address
			Heartrate_Variability_stress_level_write            => mm_interconnect_0_heartrate_variability_stress_level_write,           --                                              .write
			Heartrate_Variability_stress_level_readdata         => mm_interconnect_0_heartrate_variability_stress_level_readdata,        --                                              .readdata
			Heartrate_Variability_stress_level_writedata        => mm_interconnect_0_heartrate_variability_stress_level_writedata,       --                                              .writedata
			Interval_Timer_s1_address                           => mm_interconnect_0_interval_timer_s1_address,                          --                             Interval_Timer_s1.address
			Interval_Timer_s1_write                             => mm_interconnect_0_interval_timer_s1_write,                            --                                              .write
			Interval_Timer_s1_readdata                          => mm_interconnect_0_interval_timer_s1_readdata,                         --                                              .readdata
			Interval_Timer_s1_writedata                         => mm_interconnect_0_interval_timer_s1_writedata,                        --                                              .writedata
			Interval_Timer_s1_chipselect                        => mm_interconnect_0_interval_timer_s1_chipselect,                       --                                              .chipselect
			Interval_Timer_2_s1_address                         => mm_interconnect_0_interval_timer_2_s1_address,                        --                           Interval_Timer_2_s1.address
			Interval_Timer_2_s1_write                           => mm_interconnect_0_interval_timer_2_s1_write,                          --                                              .write
			Interval_Timer_2_s1_readdata                        => mm_interconnect_0_interval_timer_2_s1_readdata,                       --                                              .readdata
			Interval_Timer_2_s1_writedata                       => mm_interconnect_0_interval_timer_2_s1_writedata,                      --                                              .writedata
			Interval_Timer_2_s1_chipselect                      => mm_interconnect_0_interval_timer_2_s1_chipselect,                     --                                              .chipselect
			jtag_uart_0_avalon_jtag_slave_address               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,              --                 jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                --                                              .write
			jtag_uart_0_avalon_jtag_slave_read                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                 --                                              .read
			jtag_uart_0_avalon_jtag_slave_readdata              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,             --                                              .readdata
			jtag_uart_0_avalon_jtag_slave_writedata             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,            --                                              .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,          --                                              .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,           --                                              .chipselect
			nios2_gen2_0_debug_mem_slave_address                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,               --                  nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                  => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                 --                                              .write
			nios2_gen2_0_debug_mem_slave_read                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                  --                                              .read
			nios2_gen2_0_debug_mem_slave_readdata               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,              --                                              .readdata
			nios2_gen2_0_debug_mem_slave_writedata              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,             --                                              .writedata
			nios2_gen2_0_debug_mem_slave_byteenable             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,            --                                              .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,           --                                              .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,           --                                              .debugaccess
			ps2_0_avalon_ps2_slave_address                      => mm_interconnect_0_ps2_0_avalon_ps2_slave_address,                     --                        ps2_0_avalon_ps2_slave.address
			ps2_0_avalon_ps2_slave_write                        => mm_interconnect_0_ps2_0_avalon_ps2_slave_write,                       --                                              .write
			ps2_0_avalon_ps2_slave_read                         => mm_interconnect_0_ps2_0_avalon_ps2_slave_read,                        --                                              .read
			ps2_0_avalon_ps2_slave_readdata                     => mm_interconnect_0_ps2_0_avalon_ps2_slave_readdata,                    --                                              .readdata
			ps2_0_avalon_ps2_slave_writedata                    => mm_interconnect_0_ps2_0_avalon_ps2_slave_writedata,                   --                                              .writedata
			ps2_0_avalon_ps2_slave_byteenable                   => mm_interconnect_0_ps2_0_avalon_ps2_slave_byteenable,                  --                                              .byteenable
			ps2_0_avalon_ps2_slave_waitrequest                  => mm_interconnect_0_ps2_0_avalon_ps2_slave_waitrequest,                 --                                              .waitrequest
			ps2_0_avalon_ps2_slave_chipselect                   => mm_interconnect_0_ps2_0_avalon_ps2_slave_chipselect,                  --                                              .chipselect
			pushbuttons_s1_address                              => mm_interconnect_0_pushbuttons_s1_address,                             --                                pushbuttons_s1.address
			pushbuttons_s1_write                                => mm_interconnect_0_pushbuttons_s1_write,                               --                                              .write
			pushbuttons_s1_readdata                             => mm_interconnect_0_pushbuttons_s1_readdata,                            --                                              .readdata
			pushbuttons_s1_writedata                            => mm_interconnect_0_pushbuttons_s1_writedata,                           --                                              .writedata
			pushbuttons_s1_chipselect                           => mm_interconnect_0_pushbuttons_s1_chipselect,                          --                                              .chipselect
			sdram_controller_s1_address                         => mm_interconnect_0_sdram_controller_s1_address,                        --                           sdram_controller_s1.address
			sdram_controller_s1_write                           => mm_interconnect_0_sdram_controller_s1_write,                          --                                              .write
			sdram_controller_s1_read                            => mm_interconnect_0_sdram_controller_s1_read,                           --                                              .read
			sdram_controller_s1_readdata                        => mm_interconnect_0_sdram_controller_s1_readdata,                       --                                              .readdata
			sdram_controller_s1_writedata                       => mm_interconnect_0_sdram_controller_s1_writedata,                      --                                              .writedata
			sdram_controller_s1_byteenable                      => mm_interconnect_0_sdram_controller_s1_byteenable,                     --                                              .byteenable
			sdram_controller_s1_readdatavalid                   => mm_interconnect_0_sdram_controller_s1_readdatavalid,                  --                                              .readdatavalid
			sdram_controller_s1_waitrequest                     => mm_interconnect_0_sdram_controller_s1_waitrequest,                    --                                              .waitrequest
			sdram_controller_s1_chipselect                      => mm_interconnect_0_sdram_controller_s1_chipselect,                     --                                              .chipselect
			spi_0_spi_control_port_address                      => mm_interconnect_0_spi_0_spi_control_port_address,                     --                        spi_0_spi_control_port.address
			spi_0_spi_control_port_write                        => mm_interconnect_0_spi_0_spi_control_port_write,                       --                                              .write
			spi_0_spi_control_port_read                         => mm_interconnect_0_spi_0_spi_control_port_read,                        --                                              .read
			spi_0_spi_control_port_readdata                     => mm_interconnect_0_spi_0_spi_control_port_readdata,                    --                                              .readdata
			spi_0_spi_control_port_writedata                    => mm_interconnect_0_spi_0_spi_control_port_writedata,                   --                                              .writedata
			spi_0_spi_control_port_chipselect                   => mm_interconnect_0_spi_0_spi_control_port_chipselect,                  --                                              .chipselect
			spi_pio_s1_address                                  => mm_interconnect_0_spi_pio_s1_address,                                 --                                    spi_pio_s1.address
			spi_pio_s1_write                                    => mm_interconnect_0_spi_pio_s1_write,                                   --                                              .write
			spi_pio_s1_readdata                                 => mm_interconnect_0_spi_pio_s1_readdata,                                --                                              .readdata
			spi_pio_s1_writedata                                => mm_interconnect_0_spi_pio_s1_writedata,                               --                                              .writedata
			spi_pio_s1_chipselect                               => mm_interconnect_0_spi_pio_s1_chipselect,                              --                                              .chipselect
			sram_0_avalon_sram_slave_address                    => mm_interconnect_0_sram_0_avalon_sram_slave_address,                   --                      sram_0_avalon_sram_slave.address
			sram_0_avalon_sram_slave_write                      => mm_interconnect_0_sram_0_avalon_sram_slave_write,                     --                                              .write
			sram_0_avalon_sram_slave_read                       => mm_interconnect_0_sram_0_avalon_sram_slave_read,                      --                                              .read
			sram_0_avalon_sram_slave_readdata                   => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,                  --                                              .readdata
			sram_0_avalon_sram_slave_writedata                  => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,                 --                                              .writedata
			sram_0_avalon_sram_slave_byteenable                 => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,                --                                              .byteenable
			sram_0_avalon_sram_slave_readdatavalid              => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid,             --                                              .readdatavalid
			sysid_qsys_0_control_slave_address                  => mm_interconnect_0_sysid_qsys_0_control_slave_address,                 --                    sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                 => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,                --                                              .readdata
			vga_subsystem_char_buffer_control_slave_address     => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address,    --       vga_subsystem_char_buffer_control_slave.address
			vga_subsystem_char_buffer_control_slave_write       => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write,      --                                              .write
			vga_subsystem_char_buffer_control_slave_read        => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read,       --                                              .read
			vga_subsystem_char_buffer_control_slave_readdata    => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata,   --                                              .readdata
			vga_subsystem_char_buffer_control_slave_writedata   => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata,  --                                              .writedata
			vga_subsystem_char_buffer_control_slave_byteenable  => mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable, --                                              .byteenable
			vga_subsystem_char_buffer_slave_address             => mm_interconnect_0_vga_subsystem_char_buffer_slave_address,            --               vga_subsystem_char_buffer_slave.address
			vga_subsystem_char_buffer_slave_write               => mm_interconnect_0_vga_subsystem_char_buffer_slave_write,              --                                              .write
			vga_subsystem_char_buffer_slave_readdata            => mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata,           --                                              .readdata
			vga_subsystem_char_buffer_slave_writedata           => mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata,          --                                              .writedata
			vga_subsystem_char_buffer_slave_byteenable          => mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable,         --                                              .byteenable
			vga_subsystem_char_buffer_slave_chipselect          => mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect,         --                                              .chipselect
			vga_subsystem_char_buffer_slave_clken               => mm_interconnect_0_vga_subsystem_char_buffer_slave_clken,              --                                              .clken
			vga_subsystem_pixel_dma_control_slave_address       => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address,      --         vga_subsystem_pixel_dma_control_slave.address
			vga_subsystem_pixel_dma_control_slave_write         => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write,        --                                              .write
			vga_subsystem_pixel_dma_control_slave_read          => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read,         --                                              .read
			vga_subsystem_pixel_dma_control_slave_readdata      => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata,     --                                              .readdata
			vga_subsystem_pixel_dma_control_slave_writedata     => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata,    --                                              .writedata
			vga_subsystem_pixel_dma_control_slave_byteenable    => mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable,   --                                              .byteenable
			vga_subsystem_rgb_slave_read                        => mm_interconnect_0_vga_subsystem_rgb_slave_read,                       --                       vga_subsystem_rgb_slave.read
			vga_subsystem_rgb_slave_readdata                    => mm_interconnect_0_vga_subsystem_rgb_slave_readdata                    --                                              .readdata
		);

	irq_mapper : component Custom_qsys_irq_mapper
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	rst_controller : component custom_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => sys_sdram_pll_0_reset_source_reset,     -- reset_in1.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component custom_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_0_reset_source_reset,     -- reset_in0.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	sys_sdram_pll_0_reset_source_reset_ports_inv <= not sys_sdram_pll_0_reset_source_reset;

	video_pll_0_reset_source_reset_ports_inv <= not video_pll_0_reset_source_reset;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	mm_interconnect_0_spi_pio_s1_write_ports_inv <= not mm_interconnect_0_spi_pio_s1_write;

	mm_interconnect_0_pushbuttons_s1_write_ports_inv <= not mm_interconnect_0_pushbuttons_s1_write;

	mm_interconnect_0_interval_timer_s1_write_ports_inv <= not mm_interconnect_0_interval_timer_s1_write;

	mm_interconnect_0_interval_timer_2_s1_write_ports_inv <= not mm_interconnect_0_interval_timer_2_s1_write;

	mm_interconnect_0_spi_0_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_read;

	mm_interconnect_0_spi_0_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of Custom_qsys
