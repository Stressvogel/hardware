counter_fake_data_inst : counter_fake_data PORT MAP (
		clock	 => clock_sig,
		sset	 => sset_sig,
		q	 => q_sig
	);
