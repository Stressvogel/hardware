-- Computer_System_VGA_Subsystem.vhd

-- Generated using ACDS version 18.1 646

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Computer_System_VGA_Subsystem is
	port (
		pixel_dma_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => '0'); -- pixel_dma_control_slave.address
		pixel_dma_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --                        .byteenable
		pixel_dma_control_slave_read       : in  std_logic                     := '0';             --                        .read
		pixel_dma_control_slave_write      : in  std_logic                     := '0';             --                        .write
		pixel_dma_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                        .writedata
		pixel_dma_control_slave_readdata   : out std_logic_vector(31 downto 0);                    --                        .readdata
		rgb_slave_read                     : in  std_logic                     := '0';             --               rgb_slave.read
		rgb_slave_readdata                 : out std_logic_vector(31 downto 0);                    --                        .readdata
		sys_clk_clk                        : in  std_logic                     := '0';             --                 sys_clk.clk
		sys_reset_reset_n                  : in  std_logic                     := '0';             --               sys_reset.reset_n
		vga_CLK                            : out std_logic;                                        --                     vga.CLK
		vga_HS                             : out std_logic;                                        --                        .HS
		vga_VS                             : out std_logic;                                        --                        .VS
		vga_BLANK                          : out std_logic;                                        --                        .BLANK
		vga_SYNC                           : out std_logic;                                        --                        .SYNC
		vga_R                              : out std_logic_vector(7 downto 0);                     --                        .R
		vga_G                              : out std_logic_vector(7 downto 0);                     --                        .G
		vga_B                              : out std_logic_vector(7 downto 0);                     --                        .B
		vga_clk_clk                        : in  std_logic                     := '0';             --                 vga_clk.clk
		vga_reset_reset_n                  : in  std_logic                     := '0'              --               vga_reset.reset_n
	);
end entity Computer_System_VGA_Subsystem;

architecture rtl of Computer_System_VGA_Subsystem is
	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem is
		port (
			avalon_char_source_ready             : in  std_logic                     := 'X';             -- ready
			avalon_char_source_startofpacket     : out std_logic;                                        -- startofpacket
			avalon_char_source_endofpacket       : out std_logic;                                        -- endofpacket
			avalon_char_source_valid             : out std_logic;                                        -- valid
			avalon_char_source_data              : out std_logic_vector(39 downto 0);                    -- data
			char_buffer_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			char_buffer_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			char_buffer_control_slave_read       : in  std_logic                     := 'X';             -- read
			char_buffer_control_slave_write      : in  std_logic                     := 'X';             -- write
			char_buffer_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			char_buffer_control_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			char_buffer_slave_address            : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			char_buffer_slave_clken              : in  std_logic                     := 'X';             -- clken
			char_buffer_slave_chipselect         : in  std_logic                     := 'X';             -- chipselect
			char_buffer_slave_write              : in  std_logic                     := 'X';             -- write
			char_buffer_slave_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			char_buffer_slave_writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			char_buffer_slave_byteenable         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sys_clk_clk                          : in  std_logic                     := 'X';             -- clk
			sys_reset_reset_n                    : in  std_logic                     := 'X'              -- reset_n
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem;

	component Computer_System_VGA_Subsystem_VGA_Alpha_Blender is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			foreground_data          : in  std_logic_vector(39 downto 0) := (others => 'X'); -- data
			foreground_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			foreground_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			foreground_valid         : in  std_logic                     := 'X';             -- valid
			foreground_ready         : out std_logic;                                        -- ready
			background_data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			background_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			background_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			background_valid         : in  std_logic                     := 'X';             -- valid
			background_ready         : out std_logic;                                        -- ready
			output_ready             : in  std_logic                     := 'X';             -- ready
			output_data              : out std_logic_vector(29 downto 0);                    -- data
			output_startofpacket     : out std_logic;                                        -- startofpacket
			output_endofpacket       : out std_logic;                                        -- endofpacket
			output_valid             : out std_logic                                         -- valid
		);
	end component Computer_System_VGA_Subsystem_VGA_Alpha_Blender;

	component Computer_System_VGA_Subsystem_VGA_Controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component Computer_System_VGA_Subsystem_VGA_Controller;

	component Computer_System_VGA_Subsystem_VGA_Dual_Clock_FIFO is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component Computer_System_VGA_Subsystem_VGA_Dual_Clock_FIFO;

	component Computer_System_VGA_Subsystem_VGA_Pixel_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(15 downto 0);                    -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component Computer_System_VGA_Subsystem_VGA_Pixel_DMA;

	component Computer_System_VGA_Subsystem_VGA_Pixel_FIFO is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component Computer_System_VGA_Subsystem_VGA_Pixel_FIFO;

	component Computer_System_VGA_Subsystem_VGA_Pixel_RGB_Resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			slave_read               : in  std_logic                     := 'X';             -- read
			slave_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component Computer_System_VGA_Subsystem_VGA_Pixel_RGB_Resampler;

	component Computer_System_VGA_Subsystem_VGA_Pixel_Scaler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0);                    -- data
			stream_out_channel       : out std_logic_vector(1 downto 0)                      -- channel
		);
	end component Computer_System_VGA_Subsystem_VGA_Pixel_Scaler;

	component Computer_System_VGA_Subsystem_mm_interconnect_0 is
		port (
			Sys_Clk_clk_clk                                          : in  std_logic                     := 'X';             -- clk
			Char_Buf_Subsystem_sys_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			VGA_Pixel_DMA_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			VGA_Pixel_DMA_avalon_dma_master_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			VGA_Pixel_DMA_avalon_dma_master_waitrequest              : out std_logic;                                        -- waitrequest
			VGA_Pixel_DMA_avalon_dma_master_read                     : in  std_logic                     := 'X';             -- read
			VGA_Pixel_DMA_avalon_dma_master_readdata                 : out std_logic_vector(15 downto 0);                    -- readdata
			VGA_Pixel_DMA_avalon_dma_master_readdatavalid            : out std_logic;                                        -- readdatavalid
			VGA_Pixel_DMA_avalon_dma_master_lock                     : in  std_logic                     := 'X';             -- lock
			Char_Buf_Subsystem_char_buffer_control_slave_address     : out std_logic_vector(1 downto 0);                     -- address
			Char_Buf_Subsystem_char_buffer_control_slave_write       : out std_logic;                                        -- write
			Char_Buf_Subsystem_char_buffer_control_slave_read        : out std_logic;                                        -- read
			Char_Buf_Subsystem_char_buffer_control_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Char_Buf_Subsystem_char_buffer_control_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			Char_Buf_Subsystem_char_buffer_control_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			Char_Buf_Subsystem_char_buffer_slave_address             : out std_logic_vector(10 downto 0);                    -- address
			Char_Buf_Subsystem_char_buffer_slave_write               : out std_logic;                                        -- write
			Char_Buf_Subsystem_char_buffer_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Char_Buf_Subsystem_char_buffer_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			Char_Buf_Subsystem_char_buffer_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			Char_Buf_Subsystem_char_buffer_slave_chipselect          : out std_logic;                                        -- chipselect
			Char_Buf_Subsystem_char_buffer_slave_clken               : out std_logic                                         -- clken
		);
	end component Computer_System_VGA_Subsystem_mm_interconnect_0;

	component Computer_System_VGA_Subsystem_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_channel        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			out_0_data          : out std_logic_vector(29 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Computer_System_VGA_Subsystem_avalon_st_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal vga_alpha_blender_avalon_blended_source_valid                             : std_logic;                     -- VGA_Alpha_Blender:output_valid -> VGA_Dual_Clock_FIFO:stream_in_valid
	signal vga_alpha_blender_avalon_blended_source_data                              : std_logic_vector(29 downto 0); -- VGA_Alpha_Blender:output_data -> VGA_Dual_Clock_FIFO:stream_in_data
	signal vga_alpha_blender_avalon_blended_source_ready                             : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_in_ready -> VGA_Alpha_Blender:output_ready
	signal vga_alpha_blender_avalon_blended_source_startofpacket                     : std_logic;                     -- VGA_Alpha_Blender:output_startofpacket -> VGA_Dual_Clock_FIFO:stream_in_startofpacket
	signal vga_alpha_blender_avalon_blended_source_endofpacket                       : std_logic;                     -- VGA_Alpha_Blender:output_endofpacket -> VGA_Dual_Clock_FIFO:stream_in_endofpacket
	signal char_buf_subsystem_avalon_char_source_valid                               : std_logic;                     -- Char_Buf_Subsystem:avalon_char_source_valid -> VGA_Alpha_Blender:foreground_valid
	signal char_buf_subsystem_avalon_char_source_data                                : std_logic_vector(39 downto 0); -- Char_Buf_Subsystem:avalon_char_source_data -> VGA_Alpha_Blender:foreground_data
	signal char_buf_subsystem_avalon_char_source_ready                               : std_logic;                     -- VGA_Alpha_Blender:foreground_ready -> Char_Buf_Subsystem:avalon_char_source_ready
	signal char_buf_subsystem_avalon_char_source_startofpacket                       : std_logic;                     -- Char_Buf_Subsystem:avalon_char_source_startofpacket -> VGA_Alpha_Blender:foreground_startofpacket
	signal char_buf_subsystem_avalon_char_source_endofpacket                         : std_logic;                     -- Char_Buf_Subsystem:avalon_char_source_endofpacket -> VGA_Alpha_Blender:foreground_endofpacket
	signal vga_pixel_fifo_avalon_dc_buffer_source_valid                              : std_logic;                     -- VGA_Pixel_FIFO:stream_out_valid -> VGA_Pixel_RGB_Resampler:stream_in_valid
	signal vga_pixel_fifo_avalon_dc_buffer_source_data                               : std_logic_vector(15 downto 0); -- VGA_Pixel_FIFO:stream_out_data -> VGA_Pixel_RGB_Resampler:stream_in_data
	signal vga_pixel_fifo_avalon_dc_buffer_source_ready                              : std_logic;                     -- VGA_Pixel_RGB_Resampler:stream_in_ready -> VGA_Pixel_FIFO:stream_out_ready
	signal vga_pixel_fifo_avalon_dc_buffer_source_startofpacket                      : std_logic;                     -- VGA_Pixel_FIFO:stream_out_startofpacket -> VGA_Pixel_RGB_Resampler:stream_in_startofpacket
	signal vga_pixel_fifo_avalon_dc_buffer_source_endofpacket                        : std_logic;                     -- VGA_Pixel_FIFO:stream_out_endofpacket -> VGA_Pixel_RGB_Resampler:stream_in_endofpacket
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_valid                         : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_data                          : std_logic_vector(29 downto 0); -- VGA_Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_ready                         : std_logic;                     -- VGA_Controller:ready -> VGA_Dual_Clock_FIFO:stream_out_ready
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket                 : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	signal vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket                   : std_logic;                     -- VGA_Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	signal vga_pixel_dma_avalon_pixel_source_valid                                   : std_logic;                     -- VGA_Pixel_DMA:stream_valid -> VGA_Pixel_FIFO:stream_in_valid
	signal vga_pixel_dma_avalon_pixel_source_data                                    : std_logic_vector(15 downto 0); -- VGA_Pixel_DMA:stream_data -> VGA_Pixel_FIFO:stream_in_data
	signal vga_pixel_dma_avalon_pixel_source_ready                                   : std_logic;                     -- VGA_Pixel_FIFO:stream_in_ready -> VGA_Pixel_DMA:stream_ready
	signal vga_pixel_dma_avalon_pixel_source_startofpacket                           : std_logic;                     -- VGA_Pixel_DMA:stream_startofpacket -> VGA_Pixel_FIFO:stream_in_startofpacket
	signal vga_pixel_dma_avalon_pixel_source_endofpacket                             : std_logic;                     -- VGA_Pixel_DMA:stream_endofpacket -> VGA_Pixel_FIFO:stream_in_endofpacket
	signal vga_pixel_rgb_resampler_avalon_rgb_source_valid                           : std_logic;                     -- VGA_Pixel_RGB_Resampler:stream_out_valid -> VGA_Pixel_Scaler:stream_in_valid
	signal vga_pixel_rgb_resampler_avalon_rgb_source_data                            : std_logic_vector(29 downto 0); -- VGA_Pixel_RGB_Resampler:stream_out_data -> VGA_Pixel_Scaler:stream_in_data
	signal vga_pixel_rgb_resampler_avalon_rgb_source_ready                           : std_logic;                     -- VGA_Pixel_Scaler:stream_in_ready -> VGA_Pixel_RGB_Resampler:stream_out_ready
	signal vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket                   : std_logic;                     -- VGA_Pixel_RGB_Resampler:stream_out_startofpacket -> VGA_Pixel_Scaler:stream_in_startofpacket
	signal vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket                     : std_logic;                     -- VGA_Pixel_RGB_Resampler:stream_out_endofpacket -> VGA_Pixel_Scaler:stream_in_endofpacket
	signal vga_pixel_dma_avalon_dma_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:VGA_Pixel_DMA_avalon_dma_master_waitrequest -> VGA_Pixel_DMA:master_waitrequest
	signal vga_pixel_dma_avalon_dma_master_readdata                                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:VGA_Pixel_DMA_avalon_dma_master_readdata -> VGA_Pixel_DMA:master_readdata
	signal vga_pixel_dma_avalon_dma_master_address                                   : std_logic_vector(31 downto 0); -- VGA_Pixel_DMA:master_address -> mm_interconnect_0:VGA_Pixel_DMA_avalon_dma_master_address
	signal vga_pixel_dma_avalon_dma_master_read                                      : std_logic;                     -- VGA_Pixel_DMA:master_read -> mm_interconnect_0:VGA_Pixel_DMA_avalon_dma_master_read
	signal vga_pixel_dma_avalon_dma_master_readdatavalid                             : std_logic;                     -- mm_interconnect_0:VGA_Pixel_DMA_avalon_dma_master_readdatavalid -> VGA_Pixel_DMA:master_readdatavalid
	signal vga_pixel_dma_avalon_dma_master_lock                                      : std_logic;                     -- VGA_Pixel_DMA:master_arbiterlock -> mm_interconnect_0:VGA_Pixel_DMA_avalon_dma_master_lock
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_readdata   : std_logic_vector(31 downto 0); -- Char_Buf_Subsystem:char_buffer_control_slave_readdata -> mm_interconnect_0:Char_Buf_Subsystem_char_buffer_control_slave_readdata
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_control_slave_address -> Char_Buf_Subsystem:char_buffer_control_slave_address
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_read       : std_logic;                     -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_control_slave_read -> Char_Buf_Subsystem:char_buffer_control_slave_read
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_control_slave_byteenable -> Char_Buf_Subsystem:char_buffer_control_slave_byteenable
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_write      : std_logic;                     -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_control_slave_write -> Char_Buf_Subsystem:char_buffer_control_slave_write
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_control_slave_writedata -> Char_Buf_Subsystem:char_buffer_control_slave_writedata
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_slave_chipselect         : std_logic;                     -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_slave_chipselect -> Char_Buf_Subsystem:char_buffer_slave_chipselect
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_slave_readdata           : std_logic_vector(31 downto 0); -- Char_Buf_Subsystem:char_buffer_slave_readdata -> mm_interconnect_0:Char_Buf_Subsystem_char_buffer_slave_readdata
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_slave_address            : std_logic_vector(10 downto 0); -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_slave_address -> Char_Buf_Subsystem:char_buffer_slave_address
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_slave_byteenable -> Char_Buf_Subsystem:char_buffer_slave_byteenable
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_slave_write              : std_logic;                     -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_slave_write -> Char_Buf_Subsystem:char_buffer_slave_write
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_slave_writedata -> Char_Buf_Subsystem:char_buffer_slave_writedata
	signal mm_interconnect_0_char_buf_subsystem_char_buffer_slave_clken              : std_logic;                     -- mm_interconnect_0:Char_Buf_Subsystem_char_buffer_slave_clken -> Char_Buf_Subsystem:char_buffer_slave_clken
	signal vga_pixel_scaler_avalon_scaler_source_valid                               : std_logic;                     -- VGA_Pixel_Scaler:stream_out_valid -> avalon_st_adapter:in_0_valid
	signal vga_pixel_scaler_avalon_scaler_source_data                                : std_logic_vector(29 downto 0); -- VGA_Pixel_Scaler:stream_out_data -> avalon_st_adapter:in_0_data
	signal vga_pixel_scaler_avalon_scaler_source_ready                               : std_logic;                     -- avalon_st_adapter:in_0_ready -> VGA_Pixel_Scaler:stream_out_ready
	signal vga_pixel_scaler_avalon_scaler_source_channel                             : std_logic_vector(1 downto 0);  -- VGA_Pixel_Scaler:stream_out_channel -> avalon_st_adapter:in_0_channel
	signal vga_pixel_scaler_avalon_scaler_source_startofpacket                       : std_logic;                     -- VGA_Pixel_Scaler:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal vga_pixel_scaler_avalon_scaler_source_endofpacket                         : std_logic;                     -- VGA_Pixel_Scaler:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal avalon_st_adapter_out_0_valid                                             : std_logic;                     -- avalon_st_adapter:out_0_valid -> VGA_Alpha_Blender:background_valid
	signal avalon_st_adapter_out_0_data                                              : std_logic_vector(29 downto 0); -- avalon_st_adapter:out_0_data -> VGA_Alpha_Blender:background_data
	signal avalon_st_adapter_out_0_ready                                             : std_logic;                     -- VGA_Alpha_Blender:background_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                                     : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> VGA_Alpha_Blender:background_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                                       : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> VGA_Alpha_Blender:background_endofpacket
	signal rst_controller_reset_out_reset                                            : std_logic;                     -- rst_controller:reset_out -> [VGA_Alpha_Blender:reset, VGA_Dual_Clock_FIFO:reset_stream_in, VGA_Pixel_DMA:reset, VGA_Pixel_FIFO:reset_stream_in, VGA_Pixel_FIFO:reset_stream_out, VGA_Pixel_RGB_Resampler:reset, VGA_Pixel_Scaler:reset, avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:Char_Buf_Subsystem_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_0:VGA_Pixel_DMA_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                                        : std_logic;                     -- rst_controller_001:reset_out -> [VGA_Controller:reset, VGA_Dual_Clock_FIFO:reset_stream_out]
	signal sys_reset_reset_n_ports_inv                                               : std_logic;                     -- sys_reset_reset_n:inv -> rst_controller:reset_in0
	signal vga_reset_reset_n_ports_inv                                               : std_logic;                     -- vga_reset_reset_n:inv -> rst_controller_001:reset_in0

begin

	char_buf_subsystem : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem
		port map (
			avalon_char_source_ready             => char_buf_subsystem_avalon_char_source_ready,                               --        avalon_char_source.ready
			avalon_char_source_startofpacket     => char_buf_subsystem_avalon_char_source_startofpacket,                       --                          .startofpacket
			avalon_char_source_endofpacket       => char_buf_subsystem_avalon_char_source_endofpacket,                         --                          .endofpacket
			avalon_char_source_valid             => char_buf_subsystem_avalon_char_source_valid,                               --                          .valid
			avalon_char_source_data              => char_buf_subsystem_avalon_char_source_data,                                --                          .data
			char_buffer_control_slave_address    => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_address,    -- char_buffer_control_slave.address
			char_buffer_control_slave_byteenable => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_byteenable, --                          .byteenable
			char_buffer_control_slave_read       => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_read,       --                          .read
			char_buffer_control_slave_write      => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_write,      --                          .write
			char_buffer_control_slave_writedata  => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_writedata,  --                          .writedata
			char_buffer_control_slave_readdata   => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_readdata,   --                          .readdata
			char_buffer_slave_address            => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_address,            --         char_buffer_slave.address
			char_buffer_slave_clken              => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_clken,              --                          .clken
			char_buffer_slave_chipselect         => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_chipselect,         --                          .chipselect
			char_buffer_slave_write              => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_write,              --                          .write
			char_buffer_slave_readdata           => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_readdata,           --                          .readdata
			char_buffer_slave_writedata          => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_writedata,          --                          .writedata
			char_buffer_slave_byteenable         => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_byteenable,         --                          .byteenable
			sys_clk_clk                          => sys_clk_clk,                                                               --                   sys_clk.clk
			sys_reset_reset_n                    => sys_reset_reset_n                                                          --                 sys_reset.reset_n
		);

	vga_alpha_blender : component Computer_System_VGA_Subsystem_VGA_Alpha_Blender
		port map (
			clk                      => sys_clk_clk,                                           --                    clk.clk
			reset                    => rst_controller_reset_out_reset,                        --                  reset.reset
			foreground_data          => char_buf_subsystem_avalon_char_source_data,            -- avalon_foreground_sink.data
			foreground_startofpacket => char_buf_subsystem_avalon_char_source_startofpacket,   --                       .startofpacket
			foreground_endofpacket   => char_buf_subsystem_avalon_char_source_endofpacket,     --                       .endofpacket
			foreground_valid         => char_buf_subsystem_avalon_char_source_valid,           --                       .valid
			foreground_ready         => char_buf_subsystem_avalon_char_source_ready,           --                       .ready
			background_data          => avalon_st_adapter_out_0_data,                          -- avalon_background_sink.data
			background_startofpacket => avalon_st_adapter_out_0_startofpacket,                 --                       .startofpacket
			background_endofpacket   => avalon_st_adapter_out_0_endofpacket,                   --                       .endofpacket
			background_valid         => avalon_st_adapter_out_0_valid,                         --                       .valid
			background_ready         => avalon_st_adapter_out_0_ready,                         --                       .ready
			output_ready             => vga_alpha_blender_avalon_blended_source_ready,         --  avalon_blended_source.ready
			output_data              => vga_alpha_blender_avalon_blended_source_data,          --                       .data
			output_startofpacket     => vga_alpha_blender_avalon_blended_source_startofpacket, --                       .startofpacket
			output_endofpacket       => vga_alpha_blender_avalon_blended_source_endofpacket,   --                       .endofpacket
			output_valid             => vga_alpha_blender_avalon_blended_source_valid          --                       .valid
		);

	vga_controller : component Computer_System_VGA_Subsystem_VGA_Controller
		port map (
			clk           => vga_clk_clk,                                               --                clk.clk
			reset         => rst_controller_001_reset_out_reset,                        --              reset.reset
			data          => vga_dual_clock_fifo_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => vga_dual_clock_fifo_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => vga_dual_clock_fifo_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_CLK,                                                   -- external_interface.export
			VGA_HS        => vga_HS,                                                    --                   .export
			VGA_VS        => vga_VS,                                                    --                   .export
			VGA_BLANK     => vga_BLANK,                                                 --                   .export
			VGA_SYNC      => vga_SYNC,                                                  --                   .export
			VGA_R         => vga_R,                                                     --                   .export
			VGA_G         => vga_G,                                                     --                   .export
			VGA_B         => vga_B                                                      --                   .export
		);

	vga_dual_clock_fifo : component Computer_System_VGA_Subsystem_VGA_Dual_Clock_FIFO
		port map (
			clk_stream_in            => sys_clk_clk,                                               --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                            --         reset_stream_in.reset
			clk_stream_out           => vga_clk_clk,                                               --        clock_stream_out.clk
			reset_stream_out         => rst_controller_001_reset_out_reset,                        --        reset_stream_out.reset
			stream_in_ready          => vga_alpha_blender_avalon_blended_source_ready,             --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => vga_alpha_blender_avalon_blended_source_startofpacket,     --                        .startofpacket
			stream_in_endofpacket    => vga_alpha_blender_avalon_blended_source_endofpacket,       --                        .endofpacket
			stream_in_valid          => vga_alpha_blender_avalon_blended_source_valid,             --                        .valid
			stream_in_data           => vga_alpha_blender_avalon_blended_source_data,              --                        .data
			stream_out_ready         => vga_dual_clock_fifo_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => vga_dual_clock_fifo_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => vga_dual_clock_fifo_avalon_dc_buffer_source_data           --                        .data
		);

	vga_pixel_dma : component Computer_System_VGA_Subsystem_VGA_Pixel_DMA
		port map (
			clk                  => sys_clk_clk,                                     --                      clk.clk
			reset                => rst_controller_reset_out_reset,                  --                    reset.reset
			master_address       => vga_pixel_dma_avalon_dma_master_address,         --        avalon_dma_master.address
			master_waitrequest   => vga_pixel_dma_avalon_dma_master_waitrequest,     --                         .waitrequest
			master_arbiterlock   => vga_pixel_dma_avalon_dma_master_lock,            --                         .lock
			master_read          => vga_pixel_dma_avalon_dma_master_read,            --                         .read
			master_readdata      => vga_pixel_dma_avalon_dma_master_readdata,        --                         .readdata
			master_readdatavalid => vga_pixel_dma_avalon_dma_master_readdatavalid,   --                         .readdatavalid
			slave_address        => pixel_dma_control_slave_address,                 -- avalon_dma_control_slave.address
			slave_byteenable     => pixel_dma_control_slave_byteenable,              --                         .byteenable
			slave_read           => pixel_dma_control_slave_read,                    --                         .read
			slave_write          => pixel_dma_control_slave_write,                   --                         .write
			slave_writedata      => pixel_dma_control_slave_writedata,               --                         .writedata
			slave_readdata       => pixel_dma_control_slave_readdata,                --                         .readdata
			stream_ready         => vga_pixel_dma_avalon_pixel_source_ready,         --      avalon_pixel_source.ready
			stream_data          => vga_pixel_dma_avalon_pixel_source_data,          --                         .data
			stream_startofpacket => vga_pixel_dma_avalon_pixel_source_startofpacket, --                         .startofpacket
			stream_endofpacket   => vga_pixel_dma_avalon_pixel_source_endofpacket,   --                         .endofpacket
			stream_valid         => vga_pixel_dma_avalon_pixel_source_valid          --                         .valid
		);

	vga_pixel_fifo : component Computer_System_VGA_Subsystem_VGA_Pixel_FIFO
		port map (
			clk_stream_in            => sys_clk_clk,                                          --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                       --         reset_stream_in.reset
			clk_stream_out           => sys_clk_clk,                                          --        clock_stream_out.clk
			reset_stream_out         => rst_controller_reset_out_reset,                       --        reset_stream_out.reset
			stream_in_ready          => vga_pixel_dma_avalon_pixel_source_ready,              --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => vga_pixel_dma_avalon_pixel_source_startofpacket,      --                        .startofpacket
			stream_in_endofpacket    => vga_pixel_dma_avalon_pixel_source_endofpacket,        --                        .endofpacket
			stream_in_valid          => vga_pixel_dma_avalon_pixel_source_valid,              --                        .valid
			stream_in_data           => vga_pixel_dma_avalon_pixel_source_data,               --                        .data
			stream_out_ready         => vga_pixel_fifo_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => vga_pixel_fifo_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => vga_pixel_fifo_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => vga_pixel_fifo_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => vga_pixel_fifo_avalon_dc_buffer_source_data           --                        .data
		);

	vga_pixel_rgb_resampler : component Computer_System_VGA_Subsystem_VGA_Pixel_RGB_Resampler
		port map (
			clk                      => sys_clk_clk,                                             --               clk.clk
			reset                    => rst_controller_reset_out_reset,                          --             reset.reset
			stream_in_startofpacket  => vga_pixel_fifo_avalon_dc_buffer_source_startofpacket,    --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => vga_pixel_fifo_avalon_dc_buffer_source_endofpacket,      --                  .endofpacket
			stream_in_valid          => vga_pixel_fifo_avalon_dc_buffer_source_valid,            --                  .valid
			stream_in_ready          => vga_pixel_fifo_avalon_dc_buffer_source_ready,            --                  .ready
			stream_in_data           => vga_pixel_fifo_avalon_dc_buffer_source_data,             --                  .data
			slave_read               => rgb_slave_read,                                          --  avalon_rgb_slave.read
			slave_readdata           => rgb_slave_readdata,                                      --                  .readdata
			stream_out_ready         => vga_pixel_rgb_resampler_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => vga_pixel_rgb_resampler_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => vga_pixel_rgb_resampler_avalon_rgb_source_data           --                  .data
		);

	vga_pixel_scaler : component Computer_System_VGA_Subsystem_VGA_Pixel_Scaler
		port map (
			clk                      => sys_clk_clk,                                             --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                          --                reset.reset
			stream_in_startofpacket  => vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => vga_pixel_rgb_resampler_avalon_rgb_source_valid,         --                     .valid
			stream_in_ready          => vga_pixel_rgb_resampler_avalon_rgb_source_ready,         --                     .ready
			stream_in_data           => vga_pixel_rgb_resampler_avalon_rgb_source_data,          --                     .data
			stream_out_ready         => vga_pixel_scaler_avalon_scaler_source_ready,             -- avalon_scaler_source.ready
			stream_out_startofpacket => vga_pixel_scaler_avalon_scaler_source_startofpacket,     --                     .startofpacket
			stream_out_endofpacket   => vga_pixel_scaler_avalon_scaler_source_endofpacket,       --                     .endofpacket
			stream_out_valid         => vga_pixel_scaler_avalon_scaler_source_valid,             --                     .valid
			stream_out_data          => vga_pixel_scaler_avalon_scaler_source_data,              --                     .data
			stream_out_channel       => vga_pixel_scaler_avalon_scaler_source_channel            --                     .channel
		);

	mm_interconnect_0 : component Computer_System_VGA_Subsystem_mm_interconnect_0
		port map (
			Sys_Clk_clk_clk                                          => sys_clk_clk,                                                               --                                        Sys_Clk_clk.clk
			Char_Buf_Subsystem_sys_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                            -- Char_Buf_Subsystem_sys_reset_reset_bridge_in_reset.reset
			VGA_Pixel_DMA_reset_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                                            --          VGA_Pixel_DMA_reset_reset_bridge_in_reset.reset
			VGA_Pixel_DMA_avalon_dma_master_address                  => vga_pixel_dma_avalon_dma_master_address,                                   --                    VGA_Pixel_DMA_avalon_dma_master.address
			VGA_Pixel_DMA_avalon_dma_master_waitrequest              => vga_pixel_dma_avalon_dma_master_waitrequest,                               --                                                   .waitrequest
			VGA_Pixel_DMA_avalon_dma_master_read                     => vga_pixel_dma_avalon_dma_master_read,                                      --                                                   .read
			VGA_Pixel_DMA_avalon_dma_master_readdata                 => vga_pixel_dma_avalon_dma_master_readdata,                                  --                                                   .readdata
			VGA_Pixel_DMA_avalon_dma_master_readdatavalid            => vga_pixel_dma_avalon_dma_master_readdatavalid,                             --                                                   .readdatavalid
			VGA_Pixel_DMA_avalon_dma_master_lock                     => vga_pixel_dma_avalon_dma_master_lock,                                      --                                                   .lock
			Char_Buf_Subsystem_char_buffer_control_slave_address     => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_address,    --       Char_Buf_Subsystem_char_buffer_control_slave.address
			Char_Buf_Subsystem_char_buffer_control_slave_write       => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_write,      --                                                   .write
			Char_Buf_Subsystem_char_buffer_control_slave_read        => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_read,       --                                                   .read
			Char_Buf_Subsystem_char_buffer_control_slave_readdata    => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_readdata,   --                                                   .readdata
			Char_Buf_Subsystem_char_buffer_control_slave_writedata   => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_writedata,  --                                                   .writedata
			Char_Buf_Subsystem_char_buffer_control_slave_byteenable  => mm_interconnect_0_char_buf_subsystem_char_buffer_control_slave_byteenable, --                                                   .byteenable
			Char_Buf_Subsystem_char_buffer_slave_address             => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_address,            --               Char_Buf_Subsystem_char_buffer_slave.address
			Char_Buf_Subsystem_char_buffer_slave_write               => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_write,              --                                                   .write
			Char_Buf_Subsystem_char_buffer_slave_readdata            => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_readdata,           --                                                   .readdata
			Char_Buf_Subsystem_char_buffer_slave_writedata           => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_writedata,          --                                                   .writedata
			Char_Buf_Subsystem_char_buffer_slave_byteenable          => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_byteenable,         --                                                   .byteenable
			Char_Buf_Subsystem_char_buffer_slave_chipselect          => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_chipselect,         --                                                   .chipselect
			Char_Buf_Subsystem_char_buffer_slave_clken               => mm_interconnect_0_char_buf_subsystem_char_buffer_slave_clken               --                                                   .clken
		);

	avalon_st_adapter : component Computer_System_VGA_Subsystem_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 10,
			inUsePackets    => 1,
			inDataWidth     => 30,
			inChannelWidth  => 2,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 30,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => sys_clk_clk,                                         -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,                      -- in_rst_0.reset
			in_0_data           => vga_pixel_scaler_avalon_scaler_source_data,          --     in_0.data
			in_0_valid          => vga_pixel_scaler_avalon_scaler_source_valid,         --         .valid
			in_0_ready          => vga_pixel_scaler_avalon_scaler_source_ready,         --         .ready
			in_0_startofpacket  => vga_pixel_scaler_avalon_scaler_source_startofpacket, --         .startofpacket
			in_0_endofpacket    => vga_pixel_scaler_avalon_scaler_source_endofpacket,   --         .endofpacket
			in_0_channel        => vga_pixel_scaler_avalon_scaler_source_channel,       --         .channel
			out_0_data          => avalon_st_adapter_out_0_data,                        --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,                       --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,                       --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket,               --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket                  --         .endofpacket
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,    -- reset_in0.reset
			clk            => sys_clk_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => vga_reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => vga_clk_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

	vga_reset_reset_n_ports_inv <= not vga_reset_reset_n;

end architecture rtl; -- of Computer_System_VGA_Subsystem
